----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:05:08 04/30/2014 
-- Design Name: 
-- Module Name:    meomory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;
--USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity red_mem is
    Port ( clk : in  STD_LOGIC;
           addr : in  integer range 0 to 2759;
           red : out  STD_LOGIC_VECTOR (7 downto 0)
			 );
end red_mem;

architecture arch of red_mem is

   --constant ADDR_WIDTH: integer:=4;
   --constant DATA_WIDTH: integer:=3;
	constant  pic_size: integer := 2759;
   signal addr_reg: integer range 0 to pic_size;
   type myMemory is array (0 to pic_size)
        of integer range 0 to 255;
   -- ROM definition
   constant ROM: myMemory:=( 
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
248,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255,
255
);


begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   red <= std_logic_vector(to_unsigned(ROM(addr_reg),8));
	
end arch;

