----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:05:08 04/30/2014 
-- Design Name: 
-- Module Name:    meomory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;
--USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity blue_mario is
    Port ( clk : in  STD_LOGIC;
           addr : in  integer range 0 to 92159;
           blue : out  STD_LOGIC_VECTOR (7 downto 0)
			 );
end blue_mario;

architecture arch of blue_mario is

   --constant ADDR_WIDTH: integer:=4;
   --constant DATA_WIDTH: integer:=3;
	constant  pic_size: integer := 92159;
   signal addr_reg: integer range 0 to pic_size;
   type myMemory is array (0 to pic_size)
        of integer range 0 to 255;
   -- ROM definition
   constant ROM: myMemory:=( 
108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 107, 101, 99, 100, 101, 103, 103, 103, 101, 111, 118, 118, 119, 114, 105, 112, 114, 97, 114, 114, 142, 233, 247, 247, 248, 246, 249, 255, 248, 136, 114, 115, 126, 122, 137, 134, 140, 121, 113, 130, 117, 115, 108, 102, 101, 108, 113, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 110, 108, 107, 107, 107, 109, 104, 108, 105, 111, 120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 124, 115, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 138, 142, 143, 142, 141, 139, 140, 143, 137, 135, 136, 132, 134, 138, 134, 144, 138, 107, 108, 87, 102, 187, 193, 184, 182, 183, 180, 181, 177, 100, 101, 102, 107, 88, 98, 99, 111, 95, 102, 141, 141, 142, 141, 138, 136, 136, 140, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 138, 139, 137, 138, 139, 136, 141, 137, 137, 140, 0, 0, 3, 3, 0, 0, 7, 0, 5, 2, 0, 1, 1, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 7, 0, 0, 132, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 254, 250, 250, 254, 255, 255, 255, 254, 249, 255, 255, 255, 255, 255, 255, 255, 198, 70, 14, 0, 0, 32, 32, 27, 26, 20, 15, 17, 27, 0, 0, 0, 2, 0, 0, 0, 0, 0, 38, 161, 211, 231, 246, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 250, 250, 255, 255, 253, 247, 255, 255, 255, 235, 50, 28, 29, 29, 28, 25, 28, 19, 28, 25, 25, 24, 20, 21, 25, 27, 26, 30, 33, 31, 32, 28, 25, 28, 38, 43, 43, 37, 28, 27, 34, 35, 36, 27, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 28, 28, 30, 28, 25, 25, 28, 28, 25, 25, 16, 26, 43, 72, 241, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 111, 110, 103, 100, 101, 103, 104, 103, 98, 101, 110, 117, 119, 117, 114, 109, 105, 108, 96, 110, 100, 128, 228, 249, 255, 255, 251, 250, 255, 243, 144, 125, 126, 127, 133, 138, 103, 106, 102, 89, 113, 106, 108, 108, 101, 100, 107, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 132, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 135, 136, 141, 142, 141, 139, 138, 139, 138, 139, 139, 138, 134, 134, 137, 137, 137, 135, 109, 114, 97, 107, 173, 174, 180, 180, 187, 183, 173, 169, 110, 109, 105, 102, 100, 111, 90, 101, 102, 98, 136, 136, 137, 139, 140, 139, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 5, 12, 17, 15, 17, 17, 18, 17, 17, 18, 18, 23, 23, 24, 21, 17, 18, 17, 17, 20, 24, 22, 23, 14, 14, 17, 15, 21, 19, 16, 15, 19, 16, 18, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 16, 18, 15, 15, 19, 19, 16, 16, 19, 18, 29, 39, 0, 0, 145, 138, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 252, 252, 255, 255, 255, 255, 249, 250, 255, 255, 255, 255, 255, 255, 248, 206, 115, 77, 42, 18, 31, 5, 9, 9, 19, 17, 10, 18, 0, 0, 0, 0, 0, 0, 0, 9, 42, 95, 212, 250, 254, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 46, 241, 253, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 111, 117, 117, 113, 110, 108, 108, 108, 107, 104, 105, 102, 102, 107, 109, 115, 118, 108, 115, 116, 130, 110, 141, 246, 255, 255, 249, 255, 255, 255, 255, 239, 241, 243, 235, 242, 212, 117, 103, 130, 132, 113, 108, 110, 108, 101, 101, 103, 105, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 144, 130, 139, 134, 135, 130, 132, 132, 140, 127, 136, 126, 134, 135, 133, 131, 132, 132, 136, 133, 127, 135, 128, 139, 128, 132, 135, 131, 131, 128, 130, 135, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 133, 134, 138, 138, 135, 134, 132, 134, 139, 140, 133, 136, 121, 4, 0, 114, 92, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 132, 132, 134, 136, 136, 136, 136, 137, 140, 143, 142, 138, 136, 134, 135, 140, 141, 142, 126, 139, 139, 146, 186, 184, 181, 179, 188, 185, 179, 194, 176, 187, 185, 178, 192, 178, 110, 110, 137, 143, 134, 133, 132, 136, 144, 144, 139, 135, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 13, 221, 235, 241, 239, 239, 236, 235, 237, 244, 233, 242, 234, 240, 243, 240, 240, 239, 241, 243, 242, 235, 244, 232, 243, 231, 238, 241, 239, 234, 233, 235, 240, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 234, 233, 234, 236, 235, 235, 236, 235, 233, 234, 231, 226, 238, 200, 33, 0, 150, 140, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 252, 254, 255, 255, 255, 255, 255, 255, 255, 247, 213, 204, 173, 126, 90, 35, 3, 0, 19, 25, 24, 38, 11, 26, 39, 37, 45, 42, 0, 42, 143, 205, 239, 255, 255, 255, 249, 246, 253, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 115, 93, 103, 97, 92, 86, 91, 92, 97, 81, 80, 70, 80, 82, 76, 73, 71, 74, 79, 75, 63, 77, 85, 104, 90, 90, 81, 78, 90, 89, 83, 86, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 86, 91, 94, 87, 74, 70, 81, 90, 91, 85, 94, 93, 3, 32, 226, 238, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 114, 114, 113, 111, 108, 107, 107, 107, 109, 107, 98, 98, 108, 111, 112, 113, 113, 122, 133, 145, 124, 145, 227, 255, 255, 255, 255, 241, 234, 241, 233, 249, 255, 255, 251, 208, 114, 90, 116, 119, 110, 108, 114, 113, 107, 104, 104, 105, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 127, 107, 117, 112, 110, 110, 106, 111, 106, 95, 124, 110, 112, 110, 107, 109, 109, 107, 110, 112, 110, 124, 95, 106, 108, 116, 112, 113, 113, 114, 110, 117, 112, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 127, 119, 116, 118, 115, 117, 116, 109, 119, 121, 130, 120, 0, 0, 110, 97, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 133, 133, 134, 135, 136, 136, 137, 138, 142, 145, 141, 139, 142, 137, 131, 130, 139, 141, 131, 145, 150, 152, 173, 166, 172, 167, 184, 179, 167, 179, 178, 183, 166, 162, 190, 176, 109, 101, 132, 141, 139, 137, 132, 134, 141, 143, 140, 137, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 230, 244, 254, 249, 248, 248, 243, 248, 244, 234, 255, 252, 254, 252, 249, 252, 252, 250, 253, 255, 254, 255, 234, 244, 246, 255, 253, 253, 251, 251, 248, 255, 248, 248, 247, 248, 247, 248, 247, 248, 247, 248, 247, 248, 247, 248, 247, 248, 255, 249, 248, 251, 251, 253, 251, 238, 242, 243, 255, 219, 34, 5, 152, 150, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 255, 255, 247, 199, 182, 198, 207, 204, 207, 187, 144, 99, 48, 33, 20, 44, 44, 34, 36, 17, 26, 34, 38, 50, 55, 41, 93, 194, 243, 255, 255, 255, 255, 248, 244, 254, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 95, 66, 78, 71, 64, 64, 65, 70, 63, 45, 64, 46, 48, 44, 39, 38, 38, 36, 41, 41, 35, 56, 43, 63, 64, 66, 53, 56, 69, 73, 64, 67, 60, 60, 62, 60, 62, 60, 62, 60, 62, 60, 62, 60, 62, 60, 62, 60, 73, 65, 68, 66, 55, 57, 63, 59, 65, 70, 86, 92, 0, 25, 224, 246, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 103, 103, 104, 104, 101, 101, 101, 103, 104, 105, 100, 105, 119, 119, 108, 101, 91, 98, 115, 119, 99, 102, 134, 160, 168, 176, 161, 141, 129, 123, 120, 148, 165, 172, 150, 137, 128, 121, 116, 103, 98, 102, 117, 121, 115, 111, 108, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 31, 5, 10, 2, 5, 15, 5, 18, 13, 24, 103, 106, 114, 112, 109, 115, 115, 109, 112, 114, 106, 103, 24, 13, 10, 15, 7, 14, 6, 12, 5, 10, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 12, 6, 8, 19, 20, 3, 2, 15, 20, 20, 16, 12, 39, 0, 0, 112, 95, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 140, 140, 140, 139, 140, 140, 140, 142, 141, 143, 146, 138, 124, 114, 105, 101, 93, 94, 93, 92, 98, 83, 27, 33, 80, 98, 104, 109, 108, 95, 34, 37, 86, 116, 124, 131, 142, 139, 146, 142, 133, 131, 134, 136, 140, 140, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 16, 132, 141, 146, 138, 142, 151, 140, 153, 148, 161, 242, 247, 255, 253, 251, 255, 255, 251, 254, 255, 248, 243, 161, 149, 146, 152, 145, 152, 141, 145, 140, 143, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 135, 137, 150, 152, 139, 140, 153, 153, 148, 144, 138, 137, 17, 5, 147, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 254, 255, 255, 255, 254, 254, 255, 255, 255, 255, 214, 88, 34, 46, 56, 52, 53, 45, 31, 20, 5, 0, 0, 1, 4, 4, 0, 0, 0, 0, 0, 0, 49, 151, 218, 255, 255, 255, 253, 255, 255, 254, 252, 253, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 12, 0, 0, 0, 0, 0, 0, 1, 0, 0, 61, 57, 65, 60, 55, 59, 59, 53, 58, 60, 52, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 26, 228, 247, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 106, 100, 99, 101, 101, 100, 99, 99, 100, 106, 108, 105, 111, 119, 115, 109, 101, 116, 120, 129, 127, 119, 117, 123, 146, 165, 177, 162, 137, 129, 110, 109, 133, 165, 180, 146, 127, 148, 131, 108, 101, 93, 102, 112, 114, 113, 110, 108, 109, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 29, 6, 14, 8, 23, 30, 0, 6, 3, 13, 115, 110, 115, 107, 106, 113, 115, 104, 109, 113, 112, 113, 15, 1, 5, 7, 9, 19, 0, 7, 10, 13, 13, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 14, 14, 19, 10, 5, 13, 9, 0, 6, 11, 15, 5, 38, 0, 0, 115, 103, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 141, 141, 141, 141, 141, 142, 142, 142, 141, 137, 137, 137, 128, 114, 102, 113, 107, 106, 103, 100, 100, 99, 86, 37, 38, 68, 80, 104, 103, 105, 91, 38, 39, 61, 87, 137, 143, 138, 138, 133, 137, 136, 135, 135, 134, 138, 141, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 15, 129, 141, 146, 143, 155, 164, 128, 137, 132, 147, 249, 248, 251, 246, 243, 253, 252, 243, 245, 252, 248, 250, 146, 133, 135, 141, 141, 153, 125, 136, 138, 141, 140, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 140, 137, 143, 135, 134, 145, 142, 135, 139, 142, 144, 133, 138, 17, 6, 143, 139, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 252, 255, 255, 255, 254, 254, 254, 255, 247, 219, 145, 30, 0, 0, 2, 2, 3, 6, 12, 11, 14, 0, 5, 16, 11, 22, 12, 6, 5, 0, 0, 0, 61, 216, 255, 255, 252, 203, 203, 236, 252, 255, 255, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 7, 0, 0, 0, 0, 5, 0, 0, 0, 0, 76, 64, 65, 55, 51, 58, 60, 52, 57, 63, 62, 74, 0, 0, 0, 0, 0, 0, 0, 7, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 29, 226, 251, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 103, 101, 104, 104, 103, 101, 99, 100, 108, 113, 119, 119, 111, 109, 111, 115, 125, 118, 113, 106, 116, 125, 123, 135, 143, 155, 161, 145, 148, 126, 120, 135, 154, 173, 163, 135, 138, 114, 104, 122, 99, 109, 96, 93, 100, 102, 108, 111, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 136, 115, 118, 107, 117, 101, 28, 18, 14, 13, 119, 106, 115, 112, 115, 124, 126, 113, 114, 113, 108, 117, 15, 12, 118, 115, 114, 103, 30, 20, 19, 17, 14, 14, 16, 14, 16, 14, 16, 14, 16, 14, 16, 14, 16, 14, 16, 17, 129, 110, 36, 31, 110, 104, 29, 10, 116, 124, 115, 125, 0, 0, 114, 108, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 139, 140, 141, 142, 142, 145, 141, 134, 126, 119, 111, 104, 98, 97, 96, 108, 106, 104, 106, 101, 101, 86, 73, 52, 41, 81, 85, 96, 96, 72, 63, 41, 43, 117, 133, 134, 148, 105, 121, 139, 147, 143, 137, 135, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 16, 234, 248, 248, 239, 246, 232, 153, 145, 139, 142, 248, 240, 247, 247, 248, 255, 255, 248, 246, 247, 239, 249, 140, 139, 244, 244, 242, 232, 153, 144, 141, 139, 135, 135, 134, 135, 134, 135, 134, 135, 134, 135, 134, 135, 134, 135, 134, 135, 245, 225, 151, 150, 235, 233, 160, 141, 245, 252, 249, 227, 26, 1, 140, 140, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 254, 254, 255, 254, 252, 250, 251, 204, 106, 48, 26, 6, 0, 0, 0, 0, 6, 12, 0, 3, 0, 0, 0, 0, 2, 0, 0, 1, 0, 2, 0, 44, 208, 255, 255, 225, 105, 117, 207, 253, 255, 255, 252, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 95, 61, 64, 57, 65, 58, 0, 0, 0, 0, 69, 47, 52, 48, 47, 58, 60, 50, 51, 54, 49, 69, 0, 0, 85, 79, 71, 69, 13, 12, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 60, 0, 0, 71, 70, 6, 0, 80, 77, 68, 89, 0, 27, 217, 243, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 108, 108, 108, 106, 101, 103, 106, 121, 143, 141, 123, 115, 120, 126, 133, 121, 111, 103, 119, 129, 115, 121, 127, 148, 173, 170, 188, 165, 159, 164, 180, 185, 180, 150, 147, 117, 103, 119, 93, 110, 90, 88, 96, 102, 107, 112, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 132, 114, 117, 112, 127, 109, 18, 5, 19, 15, 124, 114, 124, 120, 112, 115, 115, 112, 120, 124, 114, 124, 15, 19, 113, 116, 123, 113, 18, 8, 15, 18, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 21, 126, 121, 25, 12, 126, 113, 14, 9, 118, 112, 115, 132, 0, 0, 121, 104, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 136, 137, 138, 139, 140, 139, 136, 138, 138, 126, 106, 94, 96, 99, 101, 102, 117, 112, 107, 110, 102, 108, 105, 88, 42, 22, 75, 77, 83, 86, 82, 60, 21, 23, 116, 141, 141, 146, 84, 106, 137, 151, 146, 137, 132, 133, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 231, 247, 249, 244, 255, 238, 144, 130, 144, 141, 254, 246, 255, 253, 245, 248, 248, 245, 253, 255, 246, 253, 141, 144, 240, 244, 252, 241, 142, 130, 138, 141, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 139, 243, 239, 141, 132, 249, 241, 145, 140, 250, 246, 251, 238, 18, 2, 146, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 252, 252, 255, 255, 246, 230, 205, 133, 18, 0, 10, 20, 0, 0, 0, 0, 9, 15, 0, 0, 0, 2, 0, 0, 15, 5, 7, 12, 21, 12, 0, 40, 209, 255, 248, 199, 43, 68, 193, 255, 255, 255, 250, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 79, 46, 51, 47, 64, 57, 0, 0, 0, 0, 70, 49, 56, 50, 42, 45, 45, 44, 52, 58, 51, 72, 0, 0, 73, 69, 71, 70, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 77, 67, 0, 0, 80, 70, 0, 0, 68, 55, 57, 88, 0, 25, 226, 243, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 111, 111, 113, 113, 114, 111, 107, 108, 116, 131, 204, 223, 247, 236, 144, 121, 119, 109, 106, 116, 116, 125, 111, 111, 128, 148, 184, 207, 180, 170, 190, 172, 190, 198, 207, 171, 153, 119, 81, 111, 105, 110, 108, 95, 105, 111, 115, 114, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 133, 116, 113, 114, 116, 115, 15, 14, 14, 15, 115, 116, 114, 113, 116, 115, 115, 116, 113, 114, 116, 115, 15, 14, 114, 115, 116, 114, 14, 12, 13, 14, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 11, 17, 112, 121, 8, 16, 109, 115, 114, 114, 108, 129, 0, 0, 117, 105, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 134, 134, 134, 134, 135, 136, 135, 135, 135, 135, 181, 181, 191, 181, 102, 91, 106, 107, 113, 116, 97, 106, 112, 113, 110, 75, 21, 16, 18, 20, 34, 9, 17, 15, 9, 22, 114, 151, 137, 155, 99, 101, 141, 144, 141, 137, 135, 135, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 237, 254, 251, 252, 253, 249, 145, 142, 142, 145, 249, 252, 251, 250, 253, 252, 252, 254, 251, 251, 252, 249, 146, 144, 247, 250, 252, 248, 143, 139, 141, 142, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 140, 148, 243, 252, 139, 149, 245, 253, 252, 253, 247, 238, 20, 4, 144, 136, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 252, 255, 255, 255, 253, 199, 150, 81, 44, 29, 0, 5, 14, 7, 0, 4, 5, 12, 0, 0, 2, 6, 14, 23, 0, 0, 9, 0, 10, 9, 0, 41, 195, 254, 224, 190, 49, 60, 208, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 80, 45, 42, 45, 53, 64, 0, 0, 0, 0, 68, 56, 51, 48, 53, 50, 48, 47, 44, 47, 54, 64, 0, 0, 70, 60, 56, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 78, 0, 0, 73, 69, 52, 50, 56, 93, 0, 21, 233, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 111, 111, 111, 111, 114, 113, 108, 110, 129, 138, 216, 238, 251, 242, 161, 126, 104, 106, 123, 147, 148, 141, 111, 108, 146, 179, 198, 192, 198, 199, 193, 215, 220, 205, 209, 186, 179, 156, 116, 116, 105, 107, 114, 102, 109, 111, 114, 111, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 133, 116, 113, 114, 116, 115, 15, 14, 14, 15, 115, 116, 114, 113, 116, 115, 115, 116, 113, 114, 116, 115, 15, 14, 114, 115, 116, 114, 14, 12, 13, 14, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 14, 13, 16, 108, 116, 10, 18, 105, 109, 115, 114, 108, 129, 0, 0, 117, 105, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 135, 135, 135, 135, 135, 135, 134, 133, 143, 134, 181, 178, 171, 164, 108, 96, 101, 100, 85, 89, 78, 88, 103, 98, 89, 61, 9, 0, 20, 25, 0, 4, 6, 0, 12, 34, 103, 141, 145, 148, 102, 103, 139, 141, 139, 137, 136, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 237, 254, 251, 252, 253, 249, 145, 142, 141, 144, 248, 252, 251, 250, 252, 252, 252, 254, 251, 252, 252, 249, 146, 145, 248, 251, 253, 249, 144, 139, 141, 142, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 148, 154, 242, 250, 142, 150, 241, 247, 252, 253, 248, 239, 21, 4, 144, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 252, 255, 255, 255, 255, 184, 99, 20, 0, 2, 0, 6, 48, 52, 10, 5, 8, 8, 0, 0, 2, 13, 15, 0, 0, 0, 0, 10, 16, 0, 0, 20, 152, 210, 189, 145, 33, 55, 203, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 80, 44, 41, 43, 51, 64, 0, 0, 0, 0, 69, 56, 51, 48, 54, 52, 48, 47, 42, 45, 54, 66, 0, 0, 65, 53, 51, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 77, 0, 0, 69, 63, 50, 46, 53, 90, 0, 19, 233, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 104, 104, 110, 110, 107, 110, 109, 132, 227, 255, 255, 255, 229, 212, 145, 150, 163, 188, 182, 167, 140, 150, 174, 211, 213, 220, 255, 255, 219, 227, 222, 220, 255, 255, 178, 134, 140, 111, 106, 99, 117, 109, 108, 105, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 136, 119, 116, 117, 119, 118, 18, 17, 17, 18, 118, 119, 117, 116, 119, 118, 118, 119, 116, 117, 119, 118, 18, 17, 117, 118, 119, 117, 17, 15, 16, 17, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 16, 107, 105, 24, 15, 114, 104, 20, 19, 118, 118, 111, 132, 0, 0, 121, 109, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 140, 137, 136, 135, 133, 124, 129, 191, 191, 173, 184, 174, 187, 143, 115, 40, 21, 18, 44, 94, 97, 31, 16, 5, 24, 138, 144, 18, 5, 0, 21, 143, 147, 35, 22, 95, 103, 106, 109, 141, 140, 141, 140, 140, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 235, 252, 249, 250, 251, 247, 143, 139, 139, 142, 247, 251, 249, 249, 251, 250, 251, 252, 249, 250, 250, 247, 144, 143, 247, 251, 252, 248, 142, 138, 140, 141, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 140, 242, 242, 155, 144, 243, 233, 148, 149, 249, 251, 249, 240, 19, 3, 144, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 250, 255, 255, 255, 249, 176, 97, 28, 15, 30, 29, 97, 156, 157, 35, 0, 0, 0, 9, 17, 0, 0, 1, 0, 59, 63, 0, 0, 0, 0, 45, 61, 29, 38, 72, 41, 8, 46, 189, 248, 255, 255, 251, 248, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 83, 49, 44, 47, 53, 66, 0, 2, 2, 0, 69, 56, 51, 48, 54, 53, 50, 49, 44, 49, 58, 69, 0, 0, 63, 50, 47, 56, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 78, 76, 0, 0, 81, 70, 0, 0, 59, 48, 42, 79, 0, 19, 220, 244, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 101, 103, 107, 108, 107, 108, 108, 132, 207, 232, 247, 255, 219, 212, 143, 162, 184, 219, 215, 194, 173, 174, 205, 224, 219, 222, 255, 255, 215, 217, 225, 217, 255, 255, 206, 166, 173, 116, 112, 99, 121, 112, 106, 104, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 135, 117, 116, 115, 119, 116, 18, 15, 17, 16, 118, 117, 117, 114, 119, 116, 118, 117, 116, 115, 119, 116, 18, 15, 117, 116, 119, 115, 17, 13, 16, 17, 17, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 16, 117, 113, 15, 5, 127, 116, 14, 11, 119, 119, 112, 133, 0, 0, 122, 110, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 140, 140, 139, 138, 135, 135, 130, 136, 178, 176, 171, 182, 172, 189, 141, 114, 18, 0, 0, 16, 63, 62, 17, 0, 0, 19, 133, 141, 12, 0, 0, 13, 144, 152, 18, 3, 94, 91, 107, 110, 139, 138, 142, 141, 140, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 235, 252, 249, 251, 251, 248, 143, 140, 139, 143, 247, 252, 250, 250, 251, 251, 250, 253, 249, 250, 250, 247, 143, 144, 247, 252, 253, 249, 142, 138, 140, 141, 138, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 139, 252, 250, 144, 132, 253, 242, 139, 138, 248, 251, 248, 239, 19, 2, 144, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 248, 252, 255, 255, 252, 199, 134, 65, 33, 44, 64, 135, 162, 156, 28, 0, 0, 0, 12, 14, 0, 0, 0, 0, 48, 56, 0, 0, 0, 0, 48, 58, 0, 0, 35, 0, 0, 41, 187, 248, 255, 255, 251, 248, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 85, 51, 44, 45, 53, 66, 0, 2, 2, 0, 66, 53, 47, 44, 53, 52, 52, 49, 44, 49, 60, 71, 0, 0, 61, 48, 44, 56, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 90, 85, 0, 0, 92, 80, 0, 0, 59, 46, 40, 79, 0, 21, 220, 242, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 111, 110, 106, 104, 108, 110, 108, 106, 115, 119, 144, 164, 214, 222, 166, 158, 104, 143, 173, 220, 225, 218, 215, 202, 206, 217, 232, 219, 216, 217, 200, 225, 221, 212, 209, 209, 219, 197, 158, 122, 119, 109, 124, 111, 105, 104, 111, 113, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 132, 113, 112, 111, 115, 112, 14, 11, 13, 12, 114, 113, 113, 110, 115, 112, 114, 113, 112, 111, 115, 112, 14, 11, 113, 112, 115, 111, 13, 9, 12, 13, 13, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 13, 14, 13, 5, 8, 114, 127, 8, 19, 120, 123, 119, 118, 111, 133, 0, 0, 122, 112, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 135, 135, 137, 139, 139, 138, 137, 138, 148, 139, 138, 140, 183, 190, 136, 137, 99, 90, 13, 4, 2, 0, 18, 12, 12, 7, 0, 0, 17, 25, 0, 4, 0, 0, 15, 19, 12, 29, 85, 100, 105, 106, 135, 137, 143, 142, 138, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 237, 255, 252, 254, 254, 251, 145, 143, 142, 146, 251, 255, 253, 253, 254, 253, 253, 255, 252, 253, 252, 249, 145, 146, 250, 254, 255, 251, 144, 140, 141, 143, 140, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 140, 139, 141, 139, 143, 243, 253, 132, 143, 246, 252, 250, 252, 248, 237, 18, 1, 141, 133, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 247, 245, 255, 255, 255, 234, 202, 138, 75, 79, 125, 152, 70, 46, 0, 0, 0, 0, 9, 0, 0, 0, 4, 0, 0, 0, 0, 13, 12, 0, 0, 0, 0, 0, 17, 1, 0, 35, 199, 255, 254, 249, 251, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 85, 49, 41, 40, 47, 60, 0, 0, 0, 0, 60, 45, 40, 39, 47, 50, 50, 49, 42, 47, 61, 73, 0, 0, 59, 44, 42, 54, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 91, 0, 0, 84, 74, 50, 44, 48, 88, 0, 25, 233, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 111, 110, 106, 106, 110, 111, 110, 107, 102, 107, 111, 128, 187, 195, 145, 144, 107, 137, 159, 200, 213, 223, 239, 231, 208, 211, 237, 239, 215, 210, 219, 224, 229, 235, 216, 207, 222, 188, 144, 122, 119, 110, 124, 109, 105, 104, 111, 113, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 132, 113, 110, 111, 113, 112, 12, 11, 11, 12, 112, 113, 111, 110, 113, 112, 112, 113, 110, 111, 113, 112, 12, 11, 111, 112, 113, 111, 11, 9, 10, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 12, 15, 16, 103, 116, 19, 28, 112, 111, 118, 116, 110, 132, 0, 0, 124, 112, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 135, 136, 137, 138, 138, 137, 137, 138, 142, 141, 127, 132, 188, 188, 128, 128, 100, 94, 35, 20, 2, 0, 0, 0, 2, 1, 1, 0, 0, 0, 4, 2, 0, 4, 1, 0, 3, 17, 76, 108, 104, 104, 134, 137, 143, 142, 138, 135, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 237, 255, 253, 254, 255, 251, 147, 143, 143, 147, 252, 255, 254, 253, 255, 253, 253, 255, 252, 252, 252, 249, 145, 146, 250, 254, 255, 251, 144, 139, 141, 142, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 142, 150, 152, 236, 244, 144, 154, 239, 243, 251, 253, 248, 237, 18, 0, 140, 133, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 248, 247, 252, 255, 255, 251, 240, 193, 148, 134, 146, 141, 32, 0, 0, 0, 0, 3, 12, 1, 0, 0, 13, 12, 0, 0, 1, 13, 18, 24, 6, 0, 0, 0, 1, 3, 0, 42, 203, 255, 254, 249, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 85, 49, 39, 40, 45, 60, 0, 0, 0, 0, 59, 45, 38, 39, 49, 50, 50, 49, 42, 49, 61, 75, 0, 0, 59, 44, 42, 56, 0, 5, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 61, 73, 0, 0, 72, 63, 48, 43, 51, 92, 0, 27, 235, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 104, 106, 110, 111, 113, 110, 103, 107, 106, 109, 140, 139, 108, 113, 117, 131, 141, 173, 198, 222, 230, 231, 236, 223, 224, 228, 229, 231, 223, 213, 225, 222, 222, 226, 225, 191, 154, 109, 112, 103, 119, 108, 103, 102, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 108, 111, 111, 108, 107, 106, 106, 109, 104, 106, 105, 111, 123, 0, 0, 135, 117, 114, 115, 117, 116, 16, 15, 15, 16, 116, 117, 115, 114, 117, 116, 116, 117, 114, 115, 117, 116, 16, 15, 115, 116, 117, 115, 15, 13, 14, 15, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 14, 109, 104, 18, 11, 118, 109, 20, 15, 115, 114, 108, 130, 0, 0, 125, 113, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 138, 136, 136, 136, 137, 139, 148, 146, 140, 154, 140, 102, 104, 109, 106, 84, 65, 23, 4, 0, 0, 10, 0, 0, 0, 4, 8, 0, 0, 0, 0, 4, 11, 0, 14, 91, 103, 104, 104, 137, 139, 143, 142, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 138, 139, 136, 141, 137, 137, 140, 0, 17, 235, 252, 251, 252, 253, 249, 144, 140, 140, 144, 249, 253, 252, 250, 252, 250, 251, 252, 250, 250, 250, 246, 143, 143, 248, 252, 254, 248, 141, 136, 138, 140, 138, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 138, 137, 141, 246, 244, 153, 144, 249, 241, 151, 150, 251, 253, 249, 239, 19, 1, 141, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 252, 254, 255, 255, 244, 222, 219, 171, 88, 45, 11, 3, 5, 16, 4, 5, 6, 0, 0, 0, 4, 11, 2, 1, 0, 0, 0, 0, 5, 16, 10, 0, 11, 0, 5, 62, 201, 255, 255, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 248, 250, 255, 255, 251, 247, 255, 255, 255, 228, 28, 0, 87, 51, 41, 42, 47, 60, 0, 0, 0, 0, 62, 47, 42, 42, 53, 55, 52, 51, 44, 49, 63, 76, 0, 0, 61, 46, 44, 59, 0, 9, 4, 2, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 0, 72, 59, 0, 0, 75, 70, 0, 0, 53, 46, 48, 88, 0, 23, 226, 247, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 108, 110, 113, 110, 106, 101, 102, 107, 127, 128, 107, 103, 114, 126, 147, 175, 193, 220, 227, 234, 229, 230, 225, 213, 223, 227, 222, 227, 198, 187, 172, 168, 177, 148, 127, 101, 96, 92, 114, 108, 105, 104, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 110, 110, 108, 107, 106, 107, 109, 104, 106, 103, 111, 123, 0, 0, 135, 117, 114, 117, 119, 118, 18, 17, 17, 18, 118, 119, 117, 114, 117, 116, 118, 119, 116, 117, 119, 118, 18, 17, 117, 118, 119, 117, 17, 15, 16, 17, 17, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 17, 19, 14, 114, 106, 13, 5, 120, 111, 16, 10, 115, 115, 108, 132, 0, 0, 124, 112, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 139, 136, 136, 136, 137, 137, 138, 142, 142, 146, 135, 106, 96, 103, 98, 87, 67, 21, 6, 0, 0, 0, 0, 4, 0, 0, 1, 0, 11, 7, 17, 15, 13, 10, 20, 88, 108, 101, 101, 137, 140, 142, 141, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 136, 137, 138, 139, 138, 137, 139, 136, 141, 138, 137, 140, 0, 17, 235, 252, 250, 251, 252, 248, 143, 139, 139, 142, 247, 252, 251, 250, 252, 251, 250, 252, 250, 250, 250, 246, 143, 142, 247, 251, 252, 247, 140, 136, 138, 139, 138, 138, 136, 138, 136, 138, 136, 138, 136, 138, 136, 138, 136, 138, 136, 141, 252, 248, 153, 143, 253, 243, 148, 143, 251, 252, 249, 238, 18, 1, 142, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 254, 255, 255, 255, 252, 254, 255, 255, 240, 223, 215, 161, 60, 6, 0, 0, 14, 20, 1, 6, 8, 7, 0, 0, 11, 4, 3, 2, 0, 16, 25, 43, 44, 47, 56, 43, 55, 54, 61, 106, 213, 251, 255, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 254, 250, 252, 255, 255, 251, 247, 255, 255, 255, 228, 27, 0, 87, 51, 42, 42, 49, 62, 0, 4, 4, 0, 66, 51, 43, 42, 51, 52, 52, 49, 42, 47, 60, 73, 0, 0, 61, 50, 47, 61, 0, 9, 3, 2, 1, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 0, 81, 65, 0, 0, 76, 71, 0, 0, 55, 50, 48, 86, 0, 23, 224, 247, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 107, 106, 106, 107, 107, 108, 114, 109, 121, 119, 95, 93, 108, 102, 109, 150, 165, 192, 215, 210, 218, 225, 240, 221, 217, 209, 211, 228, 231, 195, 197, 159, 155, 155, 157, 149, 129, 120, 120, 117, 111, 108, 107, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 108, 108, 107, 107, 107, 107, 109, 104, 105, 103, 109, 120, 0, 0, 132, 116, 113, 115, 119, 118, 19, 18, 18, 19, 118, 119, 115, 113, 116, 115, 116, 117, 114, 115, 117, 116, 16, 15, 115, 116, 117, 115, 15, 13, 14, 17, 16, 16, 17, 16, 17, 16, 17, 16, 17, 16, 17, 16, 17, 16, 17, 14, 6, 10, 105, 116, 7, 18, 115, 122, 119, 118, 112, 134, 0, 0, 119, 106, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 140, 138, 137, 139, 138, 139, 128, 137, 134, 109, 103, 106, 94, 94, 93, 30, 8, 11, 0, 0, 0, 0, 0, 5, 5, 0, 6, 0, 8, 108, 121, 122, 122, 120, 125, 137, 142, 141, 140, 138, 138, 138, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 140, 137, 137, 138, 138, 137, 138, 139, 136, 141, 138, 138, 142, 1, 19, 237, 253, 251, 251, 252, 247, 142, 138, 137, 141, 246, 251, 251, 252, 255, 253, 252, 253, 251, 252, 252, 249, 145, 144, 248, 251, 253, 248, 142, 138, 140, 141, 139, 139, 138, 139, 138, 139, 138, 139, 138, 139, 138, 139, 138, 139, 138, 140, 141, 150, 247, 255, 141, 148, 244, 251, 249, 250, 247, 237, 17, 0, 143, 136, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 247, 248, 255, 255, 250, 252, 255, 255, 248, 193, 83, 32, 31, 11, 3, 14, 0, 0, 4, 0, 6, 7, 8, 0, 4, 4, 0, 5, 0, 27, 172, 208, 209, 211, 213, 211, 202, 200, 206, 218, 241, 252, 254, 254, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 250, 247, 247, 254, 255, 254, 254, 255, 255, 251, 249, 255, 255, 255, 227, 27, 0, 83, 49, 41, 43, 51, 66, 0, 5, 7, 0, 71, 54, 43, 39, 42, 43, 46, 47, 39, 42, 53, 64, 0, 0, 61, 52, 49, 61, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 67, 74, 0, 0, 63, 62, 55, 53, 49, 86, 0, 25, 233, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 108, 106, 106, 104, 106, 107, 111, 114, 131, 127, 98, 95, 113, 116, 106, 146, 175, 209, 231, 222, 223, 220, 220, 200, 190, 172, 159, 166, 168, 138, 145, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 131, 113, 112, 113, 117, 116, 18, 17, 17, 18, 116, 116, 114, 112, 113, 112, 115, 116, 113, 114, 116, 115, 15, 14, 114, 115, 116, 114, 14, 12, 13, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 13, 15, 17, 105, 114, 11, 22, 114, 118, 121, 121, 115, 137, 0, 0, 119, 105, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 139, 140, 138, 139, 140, 139, 135, 129, 138, 133, 111, 106, 112, 109, 97, 85, 12, 0, 8, 0, 0, 0, 0, 0, 21, 23, 10, 13, 8, 22, 125, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 141, 141, 137, 136, 137, 138, 137, 138, 139, 136, 141, 138, 138, 142, 1, 20, 238, 255, 252, 253, 252, 248, 142, 139, 138, 142, 247, 252, 252, 252, 255, 255, 253, 254, 252, 253, 253, 250, 146, 145, 249, 252, 253, 248, 143, 139, 141, 142, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 145, 151, 243, 251, 142, 149, 239, 244, 248, 248, 245, 235, 15, 0, 142, 136, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 254, 247, 248, 255, 255, 248, 250, 255, 255, 255, 191, 58, 14, 55, 65, 54, 54, 3, 0, 9, 0, 7, 9, 12, 13, 40, 43, 39, 43, 36, 71, 220, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 250, 245, 247, 255, 255, 255, 255, 255, 255, 251, 249, 255, 255, 255, 227, 27, 0, 83, 49, 42, 43, 51, 66, 0, 5, 7, 0, 73, 56, 45, 39, 42, 43, 44, 45, 37, 40, 49, 59, 0, 0, 61, 52, 51, 63, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 70, 75, 0, 0, 57, 56, 57, 55, 51, 88, 0, 28, 236, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 108, 106, 106, 104, 104, 106, 114, 116, 128, 117, 88, 90, 122, 133, 139, 158, 171, 198, 225, 224, 225, 213, 196, 181, 182, 171, 154, 152, 147, 142, 117, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 128, 110, 109, 110, 115, 114, 15, 14, 14, 15, 114, 113, 111, 109, 110, 109, 112, 113, 110, 111, 113, 112, 12, 11, 111, 112, 113, 111, 11, 9, 10, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 13, 113, 113, 28, 18, 117, 109, 26, 25, 122, 121, 117, 139, 0, 0, 121, 107, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 138, 139, 138, 139, 140, 140, 140, 136, 140, 129, 104, 104, 123, 133, 142, 112, 24, 0, 2, 0, 0, 0, 2, 28, 90, 118, 119, 128, 128, 136, 135, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 140, 136, 136, 137, 138, 137, 138, 139, 135, 141, 138, 138, 142, 1, 20, 239, 255, 253, 254, 253, 250, 144, 140, 140, 143, 249, 253, 252, 252, 255, 255, 254, 255, 253, 254, 254, 251, 148, 147, 250, 253, 254, 250, 144, 139, 142, 143, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 238, 237, 154, 144, 243, 233, 148, 148, 247, 248, 244, 234, 14, 0, 141, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 252, 252, 255, 255, 250, 248, 255, 255, 255, 205, 93, 69, 128, 161, 183, 158, 66, 19, 5, 0, 0, 6, 29, 74, 153, 196, 211, 222, 218, 232, 245, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 254, 255, 255, 255, 255, 255, 255, 253, 251, 255, 255, 255, 227, 27, 0, 85, 51, 44, 45, 53, 66, 0, 4, 4, 0, 71, 58, 49, 46, 51, 50, 48, 45, 39, 42, 51, 60, 0, 0, 61, 53, 53, 63, 0, 3, 0, 0, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 84, 77, 0, 0, 74, 61, 0, 0, 57, 53, 51, 92, 0, 34, 238, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 104, 104, 104, 106, 112, 114, 121, 112, 91, 98, 127, 138, 122, 131, 141, 160, 178, 178, 180, 168, 147, 131, 135, 125, 108, 102, 91, 93, 104, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 128, 112, 109, 111, 115, 115, 15, 14, 15, 15, 115, 115, 111, 109, 112, 111, 112, 113, 112, 111, 115, 112, 14, 11, 113, 112, 115, 111, 13, 9, 12, 13, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 126, 123, 19, 7, 128, 117, 15, 12, 119, 118, 114, 136, 0, 0, 121, 107, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 138, 139, 140, 140, 143, 138, 139, 129, 112, 115, 133, 144, 141, 115, 38, 8, 15, 11, 17, 17, 18, 43, 104, 131, 132, 140, 137, 138, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 136, 135, 137, 138, 137, 138, 139, 135, 141, 138, 138, 142, 1, 19, 238, 254, 252, 252, 253, 249, 144, 141, 140, 144, 248, 252, 252, 252, 254, 253, 254, 255, 252, 253, 253, 251, 146, 146, 249, 252, 253, 249, 143, 139, 140, 142, 140, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 247, 245, 144, 134, 253, 242, 142, 140, 249, 251, 246, 235, 15, 0, 142, 135, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 250, 250, 255, 255, 255, 221, 143, 135, 193, 228, 233, 204, 119, 69, 46, 29, 36, 50, 74, 119, 198, 241, 255, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 253, 251, 255, 255, 255, 228, 28, 0, 89, 54, 48, 49, 54, 66, 0, 2, 2, 0, 71, 58, 52, 50, 56, 53, 48, 45, 39, 43, 53, 64, 0, 0, 63, 55, 53, 65, 0, 5, 1, 0, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 90, 82, 0, 0, 91, 76, 0, 0, 53, 50, 51, 92, 0, 30, 235, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 104, 104, 103, 104, 105, 106, 113, 114, 106, 110, 121, 118, 107, 123, 146, 164, 169, 160, 161, 154, 151, 130, 125, 112, 106, 110, 106, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 132, 116, 113, 115, 119, 119, 19, 18, 20, 19, 119, 119, 115, 113, 116, 115, 116, 117, 116, 115, 119, 116, 18, 15, 117, 116, 119, 115, 17, 13, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 14, 15, 116, 124, 3, 14, 116, 117, 112, 112, 108, 130, 0, 0, 117, 103, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 139, 139, 141, 140, 138, 135, 138, 138, 133, 133, 135, 137, 143, 145, 115, 112, 124, 121, 123, 121, 123, 118, 140, 141, 131, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 136, 136, 138, 138, 138, 138, 138, 135, 141, 138, 138, 142, 1, 18, 235, 252, 250, 250, 251, 246, 142, 139, 138, 142, 246, 250, 250, 249, 251, 251, 252, 253, 250, 251, 251, 248, 144, 144, 246, 250, 251, 247, 141, 137, 138, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 135, 141, 245, 255, 134, 145, 253, 255, 254, 254, 249, 239, 20, 3, 146, 139, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 252, 252, 254, 255, 255, 248, 204, 203, 244, 255, 253, 247, 219, 210, 209, 202, 208, 212, 225, 226, 255, 255, 255, 255, 254, 253, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 254, 255, 255, 255, 252, 255, 255, 255, 228, 30, 0, 91, 56, 50, 51, 56, 68, 0, 0, 0, 0, 69, 58, 52, 51, 60, 57, 48, 45, 41, 45, 54, 66, 0, 0, 65, 55, 53, 65, 0, 7, 3, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 64, 80, 0, 0, 62, 51, 44, 48, 49, 86, 0, 16, 226, 253, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 106, 104, 104, 104, 104, 106, 104, 106, 109, 113, 115, 116, 105, 79, 95, 116, 126, 118, 109, 112, 111, 121, 100, 99, 95, 100, 114, 109, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 132, 117, 114, 117, 120, 121, 21, 20, 21, 21, 121, 120, 117, 114, 117, 116, 118, 119, 117, 117, 120, 118, 19, 17, 118, 118, 120, 117, 18, 15, 17, 18, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 24, 23, 106, 113, 14, 22, 105, 106, 112, 112, 107, 130, 0, 0, 119, 106, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 139, 139, 139, 139, 139, 139, 139, 134, 135, 138, 143, 142, 136, 133, 126, 137, 128, 132, 137, 134, 138, 137, 145, 130, 140, 135, 130, 140, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 136, 136, 138, 139, 138, 137, 138, 134, 140, 138, 138, 141, 1, 18, 235, 251, 249, 249, 250, 246, 141, 138, 138, 142, 246, 250, 250, 249, 251, 250, 251, 253, 249, 250, 250, 247, 143, 143, 245, 249, 250, 246, 140, 136, 137, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 145, 149, 235, 246, 145, 156, 245, 249, 254, 254, 249, 239, 20, 2, 144, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 255, 255, 255, 255, 255, 255, 255, 255, 241, 245, 255, 255, 244, 249, 248, 254, 255, 253, 255, 255, 255, 252, 255, 255, 254, 255, 255, 251, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 252, 255, 255, 255, 254, 255, 255, 255, 230, 30, 0, 91, 58, 51, 52, 56, 68, 0, 0, 0, 0, 66, 54, 49, 50, 58, 55, 48, 45, 42, 47, 56, 68, 0, 0, 67, 57, 53, 65, 0, 7, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 57, 71, 0, 0, 58, 45, 46, 48, 51, 88, 0, 18, 228, 253, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 106, 106, 106, 106, 106, 111, 108, 104, 104, 108, 110, 111, 105, 100, 104, 112, 113, 104, 99, 110, 111, 111, 97, 104, 103, 106, 113, 100, 96, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 131, 115, 113, 115, 117, 118, 19, 18, 20, 19, 118, 117, 115, 113, 115, 114, 116, 117, 116, 115, 119, 116, 18, 15, 117, 116, 119, 115, 17, 13, 16, 17, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 19, 119, 115, 25, 15, 120, 109, 19, 16, 116, 116, 114, 137, 0, 0, 128, 116, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 140, 139, 139, 138, 138, 141, 138, 133, 134, 140, 142, 138, 139, 149, 151, 140, 136, 132, 129, 134, 136, 139, 130, 146, 145, 139, 146, 139, 136, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 140, 137, 137, 139, 139, 138, 137, 138, 134, 140, 137, 138, 142, 1, 18, 236, 253, 250, 250, 251, 247, 142, 139, 138, 143, 248, 252, 251, 251, 254, 252, 252, 253, 249, 250, 250, 248, 144, 144, 246, 250, 251, 247, 141, 137, 138, 139, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 239, 235, 145, 138, 247, 241, 151, 148, 250, 251, 245, 234, 13, 0, 137, 130, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 252, 250, 252, 254, 255, 255, 255, 255, 255, 255, 251, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 246, 255, 255, 255, 255, 255, 250, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 254, 255, 255, 250, 248, 255, 255, 255, 255, 255, 255, 255, 228, 30, 0, 91, 56, 50, 51, 58, 69, 0, 0, 0, 0, 64, 51, 45, 44, 51, 52, 46, 45, 44, 49, 58, 68, 0, 0, 67, 57, 53, 65, 0, 7, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 80, 75, 0, 0, 78, 69, 0, 0, 55, 50, 53, 95, 0, 34, 238, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 106, 106, 106, 107, 107, 108, 110, 109, 107, 106, 108, 106, 106, 104, 91, 92, 100, 107, 108, 109, 118, 114, 111, 96, 104, 101, 99, 108, 102, 104, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 104, 105, 102, 109, 120, 0, 0, 131, 113, 112, 114, 117, 116, 18, 18, 18, 18, 116, 117, 114, 112, 113, 114, 115, 117, 114, 115, 117, 116, 16, 15, 115, 116, 117, 115, 15, 13, 14, 15, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 124, 118, 21, 11, 121, 111, 15, 10, 118, 119, 115, 139, 0, 0, 129, 117, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 140, 140, 140, 138, 137, 136, 138, 139, 137, 136, 139, 138, 136, 140, 138, 139, 134, 136, 137, 136, 139, 135, 140, 131, 146, 141, 130, 137, 139, 141, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 140, 138, 138, 139, 139, 138, 137, 138, 134, 140, 138, 138, 142, 1, 20, 237, 254, 251, 251, 251, 248, 143, 139, 139, 143, 249, 253, 252, 252, 255, 253, 253, 253, 250, 250, 251, 248, 145, 144, 246, 250, 252, 248, 142, 137, 138, 140, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 140, 246, 240, 144, 136, 251, 243, 147, 141, 249, 250, 244, 233, 13, 0, 136, 129, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 250, 247, 248, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 253, 255, 255, 255, 255, 255, 255, 255, 247, 255, 254, 246, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 250, 254, 252, 248, 248, 255, 255, 255, 255, 255, 255, 255, 227, 28, 0, 85, 51, 46, 49, 56, 68, 0, 0, 0, 0, 62, 49, 42, 41, 47, 46, 46, 47, 46, 51, 58, 68, 0, 0, 68, 59, 54, 63, 0, 5, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 86, 79, 0, 0, 81, 71, 0, 0, 57, 50, 53, 93, 0, 30, 240, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 104, 106, 106, 107, 108, 108, 110, 110, 110, 110, 108, 108, 107, 108, 106, 103, 103, 106, 110, 114, 117, 118, 115, 108, 104, 103, 106, 114, 117, 114, 113, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 116, 109, 97, 108, 104, 117, 0, 0, 133, 110, 111, 116, 113, 113, 19, 12, 19, 15, 122, 112, 121, 117, 106, 111, 112, 109, 118, 121, 111, 121, 12, 16, 118, 114, 111, 117, 13, 19, 16, 13, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 13, 13, 12, 111, 120, 3, 14, 109, 113, 113, 119, 113, 139, 0, 0, 120, 117, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 139, 140, 140, 139, 137, 136, 135, 135, 136, 136, 137, 137, 138, 138, 140, 141, 141, 141, 139, 137, 136, 135, 135, 137, 139, 139, 138, 134, 133, 135, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 141, 141, 139, 138, 139, 139, 137, 137, 145, 139, 133, 145, 134, 140, 8, 20, 240, 253, 251, 254, 248, 245, 144, 135, 142, 140, 255, 248, 255, 255, 249, 251, 249, 246, 255, 255, 246, 255, 143, 146, 251, 249, 247, 251, 142, 145, 143, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 139, 144, 148, 246, 255, 139, 150, 250, 252, 250, 255, 248, 240, 20, 3, 135, 136, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 250, 247, 248, 254, 255, 255, 255, 255, 255, 254, 255, 254, 250, 248, 248, 248, 245, 243, 241, 241, 243, 248, 254, 255, 255, 255, 255, 255, 254, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 248, 248, 252, 252, 248, 250, 255, 255, 255, 255, 255, 255, 244, 218, 29, 0, 82, 41, 38, 45, 47, 63, 0, 0, 2, 0, 70, 44, 47, 42, 37, 41, 45, 44, 53, 59, 55, 74, 0, 0, 72, 58, 49, 66, 0, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 77, 0, 0, 75, 63, 50, 51, 49, 86, 0, 12, 226, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 104, 106, 107, 108, 108, 110, 110, 111, 111, 110, 110, 110, 108, 110, 108, 108, 107, 107, 108, 113, 115, 117, 114, 107, 104, 104, 108, 114, 115, 113, 110, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 108, 106, 100, 106, 106, 118, 0, 0, 119, 110, 116, 114, 109, 106, 13, 18, 14, 15, 117, 105, 111, 110, 108, 120, 122, 111, 111, 112, 105, 116, 12, 11, 112, 113, 112, 113, 10, 12, 11, 12, 16, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 15, 9, 15, 106, 113, 6, 14, 101, 111, 117, 111, 112, 132, 0, 0, 118, 107, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 139, 140, 139, 138, 137, 135, 135, 134, 135, 137, 137, 136, 137, 138, 140, 139, 140, 140, 140, 139, 137, 136, 136, 138, 139, 138, 136, 134, 134, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 141, 141, 138, 137, 139, 139, 137, 137, 137, 137, 137, 144, 137, 142, 8, 22, 229, 253, 255, 254, 247, 239, 138, 141, 137, 140, 249, 242, 251, 250, 251, 255, 255, 248, 247, 248, 240, 250, 143, 142, 245, 248, 248, 248, 139, 139, 138, 139, 141, 141, 140, 141, 140, 141, 140, 141, 140, 141, 140, 141, 140, 141, 140, 143, 144, 153, 242, 248, 141, 148, 237, 247, 249, 242, 246, 237, 21, 6, 140, 132, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 250, 248, 250, 255, 255, 255, 255, 255, 252, 250, 255, 255, 247, 243, 247, 245, 243, 239, 236, 236, 239, 245, 254, 255, 255, 255, 255, 255, 252, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 248, 248, 254, 254, 250, 252, 255, 255, 255, 254, 252, 255, 243, 216, 27, 0, 68, 39, 41, 41, 40, 52, 0, 0, 0, 0, 67, 40, 41, 37, 39, 54, 58, 48, 49, 52, 49, 67, 0, 0, 66, 57, 50, 60, 0, 0, 0, 0, 1, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 1, 3, 0, 0, 0, 56, 67, 0, 0, 65, 61, 52, 42, 51, 82, 0, 9, 225, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 107, 107, 108, 108, 110, 110, 111, 111, 111, 111, 111, 110, 111, 111, 114, 113, 104, 103, 106, 107, 107, 106, 104, 104, 107, 108, 108, 104, 97, 97, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 103, 107, 110, 109, 114, 119, 0, 0, 129, 112, 110, 112, 114, 114, 18, 17, 9, 20, 119, 114, 117, 111, 105, 114, 116, 108, 112, 118, 114, 118, 17, 6, 109, 113, 113, 109, 16, 11, 12, 15, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 112, 107, 19, 13, 121, 114, 22, 18, 120, 119, 131, 135, 0, 0, 111, 105, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 137, 137, 136, 135, 135, 136, 137, 137, 135, 136, 137, 137, 135, 136, 140, 141, 140, 139, 139, 139, 139, 139, 137, 137, 138, 140, 144, 143, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 140, 138, 137, 138, 138, 137, 137, 132, 139, 148, 147, 146, 143, 2, 20, 239, 254, 251, 253, 252, 248, 144, 141, 132, 145, 250, 250, 255, 250, 247, 255, 254, 244, 248, 254, 250, 252, 148, 137, 242, 248, 249, 244, 146, 139, 141, 143, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 245, 238, 144, 135, 247, 240, 145, 139, 241, 242, 255, 238, 20, 5, 142, 142, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 250, 255, 255, 255, 255, 255, 255, 248, 248, 255, 255, 250, 247, 250, 250, 252, 252, 250, 250, 250, 252, 255, 255, 255, 255, 252, 252, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 252, 255, 255, 254, 255, 255, 255, 250, 252, 255, 254, 247, 215, 21, 0, 82, 44, 35, 37, 42, 55, 0, 0, 0, 0, 72, 54, 53, 45, 41, 54, 57, 50, 54, 60, 56, 67, 0, 0, 63, 58, 51, 56, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 70, 60, 0, 0, 75, 71, 0, 0, 58, 50, 76, 97, 0, 19, 224, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 108, 108, 108, 110, 110, 110, 110, 110, 110, 110, 111, 113, 115, 113, 104, 100, 104, 104, 103, 103, 101, 104, 108, 110, 106, 100, 93, 94, 104, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 112, 111, 106, 96, 110, 115, 0, 0, 145, 131, 131, 140, 130, 128, 44, 30, 38, 49, 127, 128, 136, 133, 129, 135, 137, 131, 134, 136, 128, 125, 46, 35, 137, 135, 130, 120, 46, 36, 31, 29, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 138, 133, 38, 29, 149, 139, 38, 33, 142, 141, 132, 124, 0, 0, 110, 102, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 139, 137, 136, 137, 136, 136, 136, 138, 138, 136, 136, 136, 136, 134, 135, 139, 141, 139, 139, 140, 140, 140, 139, 137, 136, 139, 141, 144, 144, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 140, 137, 136, 138, 137, 136, 137, 141, 143, 144, 135, 142, 138, 1, 19, 227, 237, 237, 245, 235, 228, 138, 122, 128, 141, 224, 230, 239, 238, 235, 241, 239, 233, 236, 238, 230, 226, 145, 133, 237, 237, 233, 222, 144, 132, 128, 126, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 240, 233, 128, 117, 240, 230, 127, 121, 233, 235, 236, 209, 28, 1, 141, 140, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 252, 255, 255, 255, 255, 255, 255, 248, 248, 255, 255, 254, 250, 252, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 254, 253, 240, 245, 216, 30, 0, 119, 87, 77, 80, 70, 76, 14, 15, 28, 32, 91, 84, 86, 84, 83, 91, 95, 89, 92, 92, 82, 84, 19, 10, 103, 93, 80, 78, 25, 24, 15, 13, 19, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 12, 105, 98, 14, 4, 109, 103, 21, 9, 93, 85, 97, 108, 0, 30, 223, 247, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 108, 108, 108, 108, 108, 108, 108, 110, 110, 111, 108, 103, 103, 107, 108, 104, 103, 101, 103, 110, 110, 106, 101, 100, 101, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 101, 103, 104, 102, 120, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 117, 110, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 138, 138, 137, 137, 138, 137, 136, 137, 138, 138, 136, 136, 136, 137, 136, 138, 140, 139, 137, 137, 139, 140, 140, 139, 135, 135, 137, 139, 138, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 139, 137, 136, 137, 137, 136, 137, 130, 135, 142, 140, 150, 136, 2, 2, 9, 15, 17, 24, 19, 21, 13, 10, 9, 11, 28, 16, 19, 18, 17, 17, 15, 15, 15, 18, 16, 30, 13, 13, 14, 16, 18, 26, 12, 11, 12, 13, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 17, 18, 17, 15, 12, 13, 16, 19, 20, 23, 26, 39, 3, 0, 138, 139, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 252, 252, 255, 255, 255, 254, 255, 255, 250, 250, 255, 255, 255, 254, 252, 252, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 247, 246, 251, 249, 255, 229, 51, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 42, 219, 239, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 106, 106, 106, 106, 106, 107, 107, 107, 107, 107, 106, 103, 104, 111, 113, 107, 103, 101, 104, 110, 110, 104, 101, 103, 104, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 109, 110, 105, 102, 109, 96, 5, 0, 0, 11, 0, 9, 1, 6, 5, 3, 12, 3, 7, 1, 2, 3, 0, 0, 0, 1, 4, 2, 0, 4, 0, 8, 6, 1, 0, 3, 0, 2, 1, 1, 2, 2, 4, 2, 4, 2, 4, 2, 4, 2, 4, 2, 4, 2, 4, 1, 0, 0, 1, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 14, 106, 110, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 137, 137, 139, 139, 138, 138, 139, 139, 137, 137, 138, 139, 139, 139, 140, 138, 135, 135, 138, 140, 140, 139, 136, 136, 138, 139, 137, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 139, 137, 136, 137, 137, 137, 137, 138, 142, 143, 139, 137, 114, 12, 0, 0, 6, 0, 9, 3, 5, 1, 0, 3, 0, 3, 1, 3, 6, 2, 0, 0, 1, 4, 3, 2, 6, 0, 6, 6, 2, 3, 5, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 4, 3, 0, 0, 0, 0, 1, 5, 12, 9, 14, 7, 0, 11, 127, 144, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 248, 248, 255, 255, 252, 252, 255, 255, 254, 252, 255, 255, 254, 252, 250, 252, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 253, 254, 254, 255, 222, 82, 44, 45, 46, 14, 7, 0, 0, 2, 11, 24, 12, 2, 0, 0, 0, 0, 2, 4, 3, 2, 0, 0, 0, 5, 17, 8, 0, 0, 0, 9, 16, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 8, 10, 12, 8, 0, 0, 0, 0, 14, 30, 44, 82, 216, 241, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 110, 108, 108, 107, 106, 104, 104, 103, 103, 103, 103, 104, 104, 106, 104, 104, 103, 101, 106, 115, 117, 108, 104, 103, 104, 110, 108, 101, 99, 101, 103, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 104, 104, 107, 108, 107, 107, 107, 107, 110, 110, 96, 100, 112, 130, 117, 130, 143, 130, 6, 0, 0, 0, 6, 1, 5, 2, 6, 4, 7, 2, 0, 0, 0, 0, 4, 7, 4, 5, 0, 1, 2, 0, 0, 0, 3, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 3, 11, 15, 11, 8, 7, 3, 0, 0, 106, 113, 130, 114, 109, 91, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 140, 139, 137, 138, 140, 140, 139, 138, 140, 140, 140, 140, 140, 141, 141, 141, 140, 137, 132, 132, 137, 140, 140, 140, 137, 138, 142, 142, 139, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 140, 137, 137, 138, 138, 137, 137, 139, 142, 133, 136, 138, 145, 120, 126, 136, 125, 4, 0, 2, 3, 5, 0, 0, 0, 7, 7, 10, 7, 2, 1, 0, 0, 5, 10, 8, 8, 1, 1, 3, 3, 4, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 13, 139, 144, 134, 118, 144, 143, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 250, 243, 245, 255, 255, 250, 252, 255, 255, 255, 254, 254, 252, 247, 245, 247, 252, 255, 255, 255, 255, 255, 254, 254, 254, 250, 248, 250, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 254, 255, 255, 255, 255, 255, 255, 255, 255, 248, 255, 255, 255, 213, 203, 216, 192, 43, 12, 0, 0, 3, 7, 13, 8, 1, 0, 1, 3, 2, 5, 7, 5, 7, 3, 0, 0, 6, 11, 5, 0, 0, 0, 11, 13, 5, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 2, 15, 16, 4, 0, 7, 7, 5, 34, 193, 224, 234, 226, 248, 244, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 110, 108, 108, 107, 106, 104, 104, 103, 103, 103, 103, 104, 104, 106, 104, 104, 103, 103, 107, 115, 115, 110, 106, 104, 106, 110, 108, 103, 100, 103, 104, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 111, 111, 108, 108, 108, 108, 110, 111, 111, 111, 113, 114, 117, 117, 118, 117, 114, 113, 113, 113, 110, 108, 106, 106, 106, 107, 108, 110, 110, 110, 110, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 107, 108, 107, 107, 107, 107, 101, 111, 104, 112, 107, 114, 123, 132, 122, 135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 105, 118, 119, 95, 92, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 140, 139, 138, 138, 140, 140, 139, 138, 140, 140, 140, 140, 140, 141, 141, 141, 139, 137, 132, 133, 136, 139, 140, 140, 138, 139, 141, 142, 139, 139, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 138, 138, 138, 138, 136, 135, 136, 138, 139, 140, 139, 139, 138, 139, 140, 140, 138, 136, 136, 136, 139, 139, 139, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 139, 138, 137, 138, 138, 137, 137, 130, 142, 139, 146, 133, 133, 131, 135, 124, 136, 0, 3, 17, 18, 19, 18, 14, 16, 16, 16, 15, 16, 18, 22, 21, 17, 16, 18, 18, 19, 17, 16, 14, 16, 20, 19, 17, 15, 14, 14, 13, 13, 12, 13, 12, 13, 12, 13, 12, 13, 12, 13, 12, 13, 13, 14, 15, 13, 7, 6, 9, 12, 12, 10, 2, 0, 148, 135, 129, 134, 135, 143, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 248, 243, 245, 255, 255, 250, 252, 255, 255, 255, 254, 252, 250, 247, 245, 247, 252, 255, 255, 255, 255, 255, 254, 252, 250, 247, 247, 248, 252, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 254, 254, 254, 255, 255, 255, 255, 254, 254, 254, 254, 254, 252, 250, 250, 250, 250, 252, 255, 255, 252, 245, 232, 225, 224, 224, 224, 224, 225, 231, 241, 252, 255, 255, 254, 252, 255, 254, 250, 250, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 255, 255, 254, 254, 255, 255, 247, 255, 255, 255, 255, 255, 238, 232, 225, 219, 41, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 37, 231, 245, 253, 255, 248, 250, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 108, 111, 111, 108, 107, 107, 107, 108, 108, 107, 106, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 111, 122, 115, 113, 95, 117, 104, 117, 110, 111, 129, 0, 0, 6, 0, 0, 0, 0, 0, 121, 115, 108, 111, 95, 96, 108, 103, 108, 119, 108, 117, 113, 104, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 108, 110, 114, 115, 116, 126, 0, 0, 147, 129, 135, 135, 134, 130, 32, 29, 30, 33, 130, 133, 131, 131, 132, 131, 132, 131, 132, 131, 30, 32, 131, 133, 134, 130, 33, 30, 33, 33, 34, 33, 34, 33, 34, 33, 32, 35, 32, 40, 27, 29, 139, 137, 32, 34, 137, 146, 136, 139, 132, 144, 0, 0, 117, 108, 107, 110, 103, 105, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 137, 138, 139, 138, 137, 137, 138, 138, 138, 139, 139, 139, 139, 138, 138, 137, 135, 136, 137, 138, 138, 139, 138, 138, 139, 139, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 137, 137, 138, 138, 137, 136, 136, 136, 137, 137, 137, 137, 137, 136, 142, 136, 141, 128, 150, 132, 136, 127, 128, 149, 0, 2, 17, 0, 0, 0, 7, 1, 136, 128, 125, 137, 135, 140, 147, 136, 137, 144, 131, 139, 133, 126, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 137, 137, 137, 137, 137, 137, 137, 137, 138, 137, 136, 136, 136, 135, 133, 140, 0, 13, 225, 232, 235, 235, 237, 233, 131, 126, 125, 130, 232, 237, 235, 236, 235, 236, 236, 236, 234, 233, 127, 131, 232, 238, 236, 232, 130, 125, 126, 126, 124, 125, 124, 125, 125, 126, 123, 127, 122, 132, 118, 123, 233, 233, 129, 130, 228, 236, 228, 236, 235, 224, 14, 0, 143, 140, 136, 139, 135, 140, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 250, 254, 255, 252, 254, 255, 255, 255, 254, 254, 252, 252, 250, 252, 254, 255, 255, 255, 255, 254, 254, 254, 252, 252, 252, 252, 254, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 252, 252, 255, 255, 255, 255, 255, 255, 254, 254, 255, 254, 255, 245, 248, 231, 253, 242, 255, 255, 244, 236, 50, 28, 39, 19, 21, 23, 31, 44, 217, 242, 255, 255, 249, 247, 255, 252, 241, 247, 245, 255, 254, 246, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 254, 254, 255, 255, 255, 255, 248, 247, 247, 229, 34, 0, 113, 79, 85, 85, 86, 92, 14, 19, 21, 15, 96, 90, 86, 84, 84, 82, 81, 82, 86, 97, 14, 14, 90, 83, 88, 96, 17, 21, 20, 20, 24, 24, 24, 24, 22, 22, 20, 26, 24, 31, 13, 9, 111, 107, 0, 4, 109, 112, 83, 81, 84, 113, 0, 30, 228, 253, 254, 255, 254, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 117, 101, 105, 103, 106, 112, 126, 115, 127, 93, 3, 0, 0, 0, 0, 0, 0, 2, 111, 130, 125, 97, 108, 98, 97, 102, 107, 115, 108, 111, 113, 110, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 16, 20, 17, 13, 11, 17, 101, 113, 15, 22, 109, 116, 118, 116, 112, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 137, 138, 138, 138, 137, 136, 136, 136, 136, 137, 137, 137, 137, 136, 140, 124, 137, 135, 137, 135, 139, 126, 146, 120, 36, 16, 15, 18, 16, 16, 17, 36, 135, 148, 140, 121, 148, 142, 138, 137, 135, 142, 134, 136, 137, 134, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 138, 142, 139, 135, 134, 142, 227, 243, 145, 154, 238, 247, 248, 252, 251, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 250, 252, 255, 255, 255, 255, 255, 255, 254, 254, 255, 255, 254, 236, 246, 244, 245, 249, 255, 250, 238, 167, 25, 0, 0, 0, 0, 0, 0, 19, 171, 230, 255, 255, 255, 249, 255, 255, 242, 245, 247, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 1, 5, 5, 0, 0, 0, 65, 73, 0, 0, 73, 71, 52, 46, 46, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 98, 108, 111, 113, 115, 122, 110, 123, 0, 0, 125, 153, 140, 147, 133, 144, 155, 133, 0, 0, 114, 118, 108, 98, 98, 107, 103, 103, 98, 94, 106, 111, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 18, 17, 17, 12, 24, 9, 28, 17, 111, 110, 18, 16, 123, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 136, 136, 136, 137, 137, 137, 137, 137, 137, 133, 144, 145, 142, 134, 136, 118, 137, 4, 39, 191, 230, 223, 233, 221, 231, 236, 202, 20, 8, 139, 142, 141, 136, 137, 143, 135, 135, 134, 131, 138, 141, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 140, 139, 139, 134, 147, 134, 154, 147, 241, 242, 147, 147, 253, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 252, 250, 248, 252, 255, 255, 255, 255, 255, 255, 254, 254, 255, 255, 251, 255, 255, 255, 255, 255, 242, 234, 50, 23, 103, 100, 79, 84, 75, 92, 107, 109, 0, 34, 219, 248, 246, 245, 255, 255, 248, 244, 248, 246, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 3, 2, 5, 0, 5, 0, 0, 0, 71, 71, 0, 0, 57, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 106, 106, 100, 98, 116, 106, 133, 121, 124, 0, 0, 124, 139, 124, 127, 118, 129, 123, 137, 0, 0, 113, 107, 123, 118, 96, 107, 108, 107, 107, 93, 97, 98, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 16, 14, 25, 7, 25, 7, 122, 117, 11, 6, 121, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 137, 136, 136, 136, 137, 137, 138, 138, 137, 138, 146, 140, 129, 141, 123, 148, 139, 154, 17, 41, 220, 251, 245, 252, 246, 252, 237, 238, 46, 33, 145, 129, 150, 149, 131, 141, 139, 140, 148, 135, 138, 135, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 139, 139, 138, 136, 148, 132, 151, 137, 252, 249, 140, 137, 251, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 248, 248, 252, 255, 255, 255, 255, 255, 254, 252, 252, 255, 255, 255, 255, 254, 255, 229, 239, 215, 192, 0, 0, 71, 61, 44, 47, 47, 58, 51, 84, 0, 4, 184, 212, 253, 255, 251, 255, 255, 255, 255, 253, 254, 250, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 2, 2, 4, 0, 6, 0, 0, 0, 82, 78, 0, 0, 55, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 100, 92, 128, 120, 0, 0, 0, 0, 153, 116, 140, 109, 108, 106, 113, 109, 111, 126, 121, 124, 0, 0, 117, 107, 111, 105, 109, 96, 100, 92, 103, 107, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 12, 20, 15, 12, 11, 18, 108, 122, 7, 12, 121, 126, 114, 115, 111, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 137, 137, 136, 136, 137, 137, 138, 138, 138, 138, 137, 133, 123, 152, 143, 6, 8, 24, 23, 233, 218, 255, 247, 253, 252, 255, 252, 251, 252, 226, 198, 32, 0, 135, 128, 140, 137, 138, 128, 141, 138, 146, 147, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 134, 142, 137, 134, 134, 143, 234, 252, 137, 144, 250, 255, 244, 251, 250, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 248, 248, 250, 254, 255, 255, 255, 255, 255, 252, 252, 252, 252, 255, 255, 250, 255, 223, 50, 19, 10, 0, 136, 74, 69, 27, 28, 29, 43, 38, 30, 56, 81, 121, 35, 64, 243, 253, 255, 250, 255, 251, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 5, 3, 0, 0, 0, 72, 82, 0, 0, 85, 81, 48, 45, 45, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 115, 111, 92, 0, 0, 0, 0, 122, 122, 111, 106, 115, 100, 112, 105, 109, 102, 140, 149, 0, 0, 129, 112, 109, 96, 132, 111, 101, 93, 96, 99, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 11, 19, 13, 14, 13, 15, 105, 112, 17, 19, 113, 117, 113, 115, 112, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 137, 137, 136, 136, 137, 137, 138, 138, 138, 138, 137, 135, 140, 134, 118, 34, 22, 38, 39, 227, 243, 249, 255, 255, 252, 255, 253, 255, 243, 255, 238, 16, 1, 142, 131, 140, 128, 156, 137, 140, 136, 139, 139, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 133, 141, 135, 136, 136, 140, 231, 242, 147, 151, 242, 248, 243, 251, 251, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 252, 252, 254, 255, 255, 255, 255, 255, 254, 252, 250, 250, 252, 255, 255, 255, 212, 151, 14, 0, 0, 0, 75, 62, 39, 29, 39, 29, 46, 35, 30, 25, 80, 120, 0, 44, 244, 249, 231, 215, 255, 255, 255, 255, 254, 250, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 4, 1, 0, 0, 0, 69, 72, 0, 0, 77, 72, 47, 45, 46, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 117, 104, 0, 0, 140, 156, 142, 126, 119, 126, 104, 112, 110, 108, 114, 113, 104, 117, 115, 122, 0, 0, 114, 126, 0, 0, 103, 113, 109, 105, 101, 101, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 13, 17, 13, 13, 25, 7, 32, 16, 114, 107, 22, 16, 118, 115, 115, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 137, 137, 137, 138, 138, 138, 138, 137, 139, 125, 10, 35, 194, 232, 239, 240, 244, 255, 245, 255, 253, 249, 250, 250, 248, 255, 246, 222, 33, 11, 130, 146, 9, 22, 127, 135, 140, 142, 137, 137, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 135, 139, 135, 135, 148, 132, 158, 146, 244, 239, 151, 147, 248, 251, 254, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 252, 250, 250, 252, 254, 255, 216, 48, 13, 108, 100, 82, 66, 62, 68, 42, 49, 47, 48, 54, 50, 36, 46, 44, 70, 0, 25, 215, 241, 57, 61, 199, 237, 255, 255, 255, 251, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 2, 1, 0, 6, 0, 0, 0, 74, 68, 0, 0, 52, 45, 49, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 111, 109, 116, 0, 0, 149, 141, 119, 115, 109, 114, 103, 120, 102, 119, 114, 119, 112, 112, 119, 137, 0, 0, 118, 110, 0, 0, 117, 121, 103, 104, 103, 113, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 15, 18, 16, 3, 27, 12, 12, 11, 116, 115, 16, 10, 121, 114, 114, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 136, 136, 136, 136, 136, 137, 137, 137, 137, 137, 137, 137, 137, 136, 129, 137, 6, 20, 221, 237, 239, 248, 247, 255, 246, 255, 243, 255, 247, 253, 250, 251, 254, 248, 32, 16, 150, 144, 16, 21, 147, 144, 128, 132, 135, 146, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 137, 140, 138, 125, 150, 137, 138, 141, 246, 247, 145, 141, 251, 250, 253, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 254, 254, 254, 255, 254, 244, 220, 23, 0, 96, 67, 45, 45, 47, 55, 44, 61, 42, 60, 58, 62, 51, 44, 38, 66, 0, 0, 189, 190, 5, 2, 173, 214, 244, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 4, 0, 8, 0, 0, 0, 76, 76, 0, 0, 55, 44, 48, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 99, 107, 112, 103, 114, 106, 105, 118, 117, 117, 0, 0, 139, 142, 108, 115, 111, 106, 114, 110, 114, 109, 116, 113, 119, 110, 118, 124, 138, 143, 0, 0, 146, 144, 0, 0, 105, 117, 102, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 14, 18, 14, 23, 9, 12, 121, 118, 13, 14, 115, 123, 115, 117, 113, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 136, 136, 136, 136, 137, 137, 128, 136, 141, 131, 142, 134, 133, 142, 135, 138, 8, 23, 224, 252, 238, 255, 253, 248, 253, 250, 255, 252, 255, 249, 254, 245, 255, 248, 228, 212, 22, 21, 220, 212, 17, 6, 129, 142, 130, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 136, 140, 136, 145, 132, 137, 247, 248, 143, 146, 244, 254, 245, 253, 252, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 246, 254, 255, 254, 255, 255, 255, 255, 255, 227, 25, 0, 95, 77, 41, 47, 47, 42, 46, 40, 46, 46, 61, 61, 66, 46, 34, 40, 79, 123, 0, 0, 135, 125, 0, 30, 215, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 2, 8, 0, 0, 85, 78, 0, 0, 79, 78, 49, 47, 47, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 110, 108, 105, 112, 105, 106, 110, 118, 120, 0, 0, 133, 120, 124, 110, 120, 111, 117, 115, 115, 113, 116, 108, 118, 110, 124, 119, 139, 128, 0, 0, 137, 139, 0, 0, 114, 126, 107, 105, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 16, 20, 17, 13, 11, 17, 101, 113, 15, 22, 109, 116, 118, 116, 112, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 136, 136, 136, 137, 137, 137, 136, 138, 136, 133, 139, 133, 134, 131, 128, 135, 12, 38, 227, 240, 255, 255, 255, 250, 254, 253, 255, 255, 255, 247, 246, 240, 255, 252, 249, 224, 46, 37, 235, 228, 35, 31, 140, 149, 133, 134, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 138, 142, 139, 135, 134, 142, 227, 243, 145, 154, 238, 247, 248, 252, 251, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 255, 255, 255, 255, 255, 255, 255, 255, 230, 24, 0, 91, 57, 57, 44, 56, 47, 50, 46, 46, 46, 62, 60, 71, 54, 46, 37, 72, 88, 0, 0, 90, 84, 0, 4, 189, 245, 252, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 1, 5, 5, 0, 0, 0, 65, 73, 0, 0, 73, 71, 52, 46, 46, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 112, 108, 99, 102, 104, 104, 112, 111, 126, 137, 0, 0, 143, 116, 113, 107, 109, 111, 124, 117, 110, 101, 111, 112, 18, 18, 108, 120, 105, 132, 119, 129, 120, 138, 146, 143, 0, 0, 105, 109, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 18, 17, 17, 12, 24, 9, 28, 17, 111, 110, 18, 16, 123, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 137, 137, 137, 137, 137, 141, 136, 126, 129, 131, 131, 140, 131, 125, 141, 8, 27, 241, 239, 253, 255, 250, 249, 255, 252, 250, 243, 254, 251, 144, 143, 246, 255, 235, 252, 233, 243, 241, 249, 231, 202, 16, 0, 133, 140, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 140, 139, 139, 134, 147, 134, 154, 147, 241, 242, 147, 147, 253, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 238, 16, 0, 96, 47, 42, 39, 47, 52, 63, 53, 40, 33, 52, 64, 0, 0, 47, 52, 41, 77, 83, 86, 48, 59, 88, 122, 17, 62, 242, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 3, 2, 5, 0, 5, 0, 0, 0, 71, 71, 0, 0, 57, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 103, 105, 102, 115, 109, 109, 111, 107, 126, 111, 0, 0, 126, 116, 115, 115, 102, 109, 112, 104, 120, 111, 109, 116, 12, 27, 105, 120, 110, 102, 128, 115, 119, 114, 137, 154, 0, 0, 122, 103, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 16, 14, 25, 7, 25, 7, 122, 117, 11, 6, 121, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 137, 131, 133, 129, 142, 136, 137, 141, 128, 129, 121, 37, 36, 228, 240, 253, 255, 243, 247, 244, 237, 255, 249, 248, 251, 136, 153, 240, 255, 250, 238, 255, 245, 254, 242, 242, 229, 18, 3, 152, 135, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 139, 139, 138, 136, 148, 132, 151, 137, 252, 249, 140, 137, 251, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 254, 252, 252, 252, 254, 254, 255, 255, 255, 255, 255, 255, 235, 234, 180, 10, 0, 66, 42, 43, 50, 51, 65, 64, 50, 52, 39, 45, 63, 0, 0, 59, 66, 53, 44, 69, 49, 37, 31, 64, 110, 0, 39, 248, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 2, 2, 4, 0, 6, 0, 0, 0, 82, 78, 0, 0, 55, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 114, 112, 104, 109, 98, 109, 106, 117, 0, 0, 130, 148, 145, 125, 124, 99, 19, 22, 11, 29, 110, 127, 115, 116, 116, 109, 19, 2, 113, 108, 115, 115, 105, 124, 126, 139, 0, 0, 108, 112, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 12, 20, 15, 12, 11, 18, 108, 122, 7, 12, 121, 126, 114, 115, 111, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 142, 139, 131, 136, 127, 139, 139, 146, 2, 28, 189, 231, 255, 252, 255, 239, 157, 158, 141, 159, 240, 255, 244, 245, 242, 237, 151, 140, 255, 248, 248, 249, 249, 255, 248, 228, 29, 5, 135, 142, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 134, 142, 137, 134, 134, 143, 234, 252, 137, 144, 250, 255, 244, 251, 250, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 250, 250, 254, 255, 255, 255, 255, 247, 249, 234, 216, 39, 10, 99, 87, 70, 47, 56, 46, 0, 0, 0, 0, 44, 52, 38, 54, 80, 80, 0, 0, 66, 51, 45, 38, 29, 48, 53, 84, 0, 21, 222, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 5, 3, 0, 0, 0, 72, 82, 0, 0, 85, 81, 48, 45, 45, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 106, 105, 104, 109, 109, 127, 94, 109, 0, 0, 132, 145, 109, 128, 112, 122, 5, 11, 0, 20, 104, 126, 114, 119, 114, 116, 17, 10, 117, 109, 122, 117, 112, 104, 117, 146, 0, 0, 125, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 11, 19, 13, 14, 13, 15, 105, 112, 17, 19, 113, 117, 113, 115, 112, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 134, 133, 131, 137, 139, 160, 130, 150, 18, 36, 220, 250, 229, 255, 246, 255, 142, 147, 134, 153, 236, 255, 241, 246, 245, 246, 145, 144, 255, 249, 252, 251, 255, 248, 248, 243, 21, 4, 150, 135, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 133, 141, 135, 136, 136, 140, 231, 242, 147, 151, 242, 248, 243, 251, 251, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 250, 250, 254, 255, 255, 255, 255, 249, 253, 206, 182, 0, 0, 74, 70, 33, 55, 53, 76, 0, 0, 0, 0, 38, 48, 38, 53, 69, 78, 0, 0, 70, 52, 42, 34, 42, 37, 46, 86, 0, 14, 234, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 4, 1, 0, 0, 0, 69, 72, 0, 0, 77, 72, 47, 45, 46, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 105, 106, 112, 111, 106, 94, 0, 0, 145, 111, 131, 115, 120, 126, 14, 5, 113, 113, 105, 100, 126, 121, 115, 117, 113, 122, 113, 120, 113, 102, 129, 116, 107, 115, 106, 133, 0, 0, 119, 118, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 13, 17, 13, 13, 25, 7, 32, 16, 114, 107, 22, 16, 118, 115, 115, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 137, 133, 134, 140, 140, 139, 130, 21, 22, 233, 224, 255, 248, 254, 255, 143, 136, 250, 254, 247, 242, 255, 255, 245, 248, 249, 255, 240, 247, 248, 233, 251, 240, 246, 255, 243, 234, 22, 7, 136, 140, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 135, 139, 135, 135, 148, 132, 158, 146, 244, 239, 151, 147, 248, 251, 254, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 252, 252, 252, 255, 255, 255, 255, 255, 234, 204, 73, 15, 129, 56, 62, 43, 59, 72, 0, 0, 76, 77, 64, 44, 52, 42, 48, 56, 53, 61, 45, 54, 58, 41, 44, 30, 43, 59, 43, 80, 0, 23, 224, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 2, 1, 0, 6, 0, 0, 0, 74, 68, 0, 0, 52, 45, 49, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 107, 107, 107, 108, 108, 107, 106, 106, 107, 110, 111, 120, 111, 114, 109, 117, 109, 0, 0, 127, 112, 108, 110, 103, 112, 20, 17, 117, 107, 111, 109, 114, 111, 118, 111, 115, 116, 118, 124, 115, 122, 127, 126, 111, 115, 112, 137, 0, 0, 122, 117, 111, 108, 108, 110, 113, 113, 110, 110, 111, 111, 107, 107, 111, 111, 107, 106, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 15, 18, 16, 3, 27, 12, 12, 11, 116, 115, 16, 10, 121, 114, 114, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 137, 137, 136, 137, 139, 139, 138, 137, 137, 138, 146, 136, 134, 131, 147, 150, 21, 31, 242, 249, 251, 254, 241, 246, 149, 148, 252, 248, 255, 252, 255, 250, 253, 245, 254, 252, 247, 252, 249, 254, 250, 249, 247, 255, 251, 249, 28, 10, 141, 136, 136, 137, 137, 138, 139, 139, 138, 136, 136, 136, 139, 139, 136, 136, 138, 139, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 137, 140, 138, 125, 150, 137, 138, 141, 246, 247, 145, 141, 251, 250, 253, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 252, 252, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 252, 254, 255, 255, 254, 245, 243, 229, 229, 216, 209, 182, 16, 0, 89, 45, 37, 42, 44, 61, 0, 0, 71, 58, 57, 46, 39, 37, 55, 50, 49, 46, 43, 53, 54, 56, 45, 44, 51, 60, 48, 79, 0, 0, 199, 238, 252, 255, 255, 247, 234, 234, 248, 255, 254, 254, 252, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 4, 0, 8, 0, 0, 0, 76, 76, 0, 0, 55, 44, 48, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 107, 107, 107, 107, 107, 106, 106, 106, 104, 104, 103, 106, 108, 112, 97, 92, 105, 109, 104, 115, 0, 0, 0, 0, 0, 0, 134, 132, 120, 114, 113, 113, 114, 114, 115, 114, 114, 113, 113, 113, 114, 114, 114, 114, 114, 115, 117, 115, 114, 114, 118, 118, 114, 120, 109, 118, 136, 159, 0, 0, 117, 107, 109, 115, 0, 0, 119, 107, 114, 115, 106, 106, 114, 111, 106, 104, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 14, 18, 14, 23, 9, 12, 121, 118, 13, 14, 115, 123, 115, 117, 113, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 140, 139, 139, 139, 138, 138, 138, 138, 139, 139, 139, 139, 138, 139, 137, 133, 138, 136, 135, 142, 138, 129, 137, 1, 6, 0, 4, 5, 18, 214, 240, 245, 251, 252, 252, 251, 250, 249, 250, 250, 251, 251, 252, 252, 252, 251, 251, 251, 250, 249, 250, 252, 252, 250, 249, 248, 255, 252, 246, 231, 222, 10, 6, 141, 136, 138, 141, 3, 0, 143, 129, 130, 134, 140, 140, 130, 130, 142, 146, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 136, 140, 136, 145, 132, 137, 247, 248, 143, 146, 244, 254, 245, 253, 252, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 248, 247, 248, 250, 252, 254, 255, 255, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 237, 240, 255, 255, 245, 222, 46, 34, 38, 37, 12, 0, 119, 95, 65, 49, 45, 47, 51, 54, 54, 56, 54, 52, 51, 49, 45, 45, 51, 51, 51, 51, 51, 49, 45, 43, 43, 47, 53, 59, 38, 47, 77, 131, 0, 62, 249, 255, 255, 236, 56, 55, 243, 251, 252, 252, 248, 250, 252, 251, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 2, 8, 0, 0, 85, 78, 0, 0, 79, 78, 49, 47, 47, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 107, 107, 107, 107, 107, 107, 106, 106, 104, 104, 104, 103, 103, 104, 117, 119, 108, 106, 98, 104, 113, 121, 0, 0, 0, 0, 0, 0, 118, 121, 115, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 115, 114, 113, 113, 113, 114, 115, 114, 118, 107, 115, 131, 150, 0, 0, 126, 109, 109, 105, 0, 0, 114, 114, 120, 115, 105, 102, 117, 118, 101, 101, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 16, 20, 17, 13, 11, 17, 101, 113, 15, 22, 109, 116, 118, 116, 112, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 140, 139, 139, 139, 138, 138, 138, 139, 139, 139, 139, 139, 139, 139, 139, 143, 146, 146, 147, 128, 131, 138, 149, 16, 16, 12, 14, 26, 58, 225, 250, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 250, 250, 252, 253, 253, 252, 250, 248, 255, 251, 253, 248, 234, 18, 4, 146, 133, 139, 138, 11, 12, 143, 136, 133, 135, 139, 135, 132, 133, 138, 143, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 138, 142, 139, 135, 134, 142, 227, 243, 145, 154, 238, 247, 248, 252, 251, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 247, 247, 248, 250, 252, 254, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 247, 253, 255, 255, 228, 189, 0, 0, 0, 0, 0, 0, 69, 61, 52, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 51, 52, 49, 42, 40, 45, 49, 55, 55, 31, 36, 58, 97, 0, 24, 243, 255, 235, 189, 0, 4, 201, 235, 245, 248, 247, 248, 255, 255, 252, 251, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 1, 5, 5, 0, 0, 0, 65, 73, 0, 0, 73, 71, 52, 46, 46, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 107, 107, 107, 107, 107, 107, 106, 106, 106, 104, 104, 103, 103, 104, 95, 100, 115, 97, 132, 122, 0, 0, 153, 147, 152, 140, 130, 98, 128, 107, 113, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 115, 114, 113, 113, 113, 114, 115, 116, 117, 107, 115, 128, 136, 0, 0, 109, 119, 0, 0, 154, 142, 0, 0, 109, 108, 114, 109, 114, 114, 99, 101, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 18, 17, 17, 12, 24, 9, 28, 17, 111, 110, 18, 16, 123, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 139, 140, 139, 139, 139, 138, 138, 138, 138, 138, 138, 139, 140, 141, 142, 141, 127, 127, 142, 119, 147, 140, 5, 17, 218, 224, 232, 228, 228, 213, 255, 252, 252, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 250, 250, 251, 253, 253, 252, 250, 247, 252, 251, 255, 248, 229, 32, 9, 125, 138, 5, 27, 220, 204, 22, 3, 131, 130, 141, 137, 131, 133, 132, 140, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 140, 139, 139, 134, 147, 134, 154, 147, 241, 242, 147, 147, 253, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 248, 250, 250, 252, 254, 255, 255, 255, 255, 255, 255, 252, 248, 243, 245, 238, 244, 255, 238, 255, 238, 41, 0, 124, 94, 99, 89, 79, 47, 73, 50, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 52, 51, 43, 42, 45, 49, 55, 53, 32, 36, 52, 76, 0, 4, 210, 240, 50, 4, 122, 107, 7, 47, 216, 239, 255, 255, 255, 255, 245, 243, 250, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 3, 2, 5, 0, 5, 0, 0, 0, 71, 71, 0, 0, 57, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 107, 107, 107, 107, 107, 107, 106, 106, 106, 106, 106, 104, 104, 104, 113, 103, 122, 111, 122, 117, 0, 0, 139, 126, 135, 121, 127, 113, 108, 105, 111, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 113, 111, 111, 113, 114, 115, 111, 118, 120, 124, 124, 112, 0, 0, 129, 103, 0, 0, 134, 161, 0, 0, 122, 104, 108, 106, 106, 114, 112, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 16, 14, 25, 7, 25, 7, 122, 117, 11, 6, 121, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 140, 139, 139, 139, 138, 138, 137, 138, 138, 138, 138, 140, 141, 143, 143, 150, 135, 144, 128, 139, 144, 28, 41, 229, 234, 252, 247, 255, 254, 255, 254, 252, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 253, 252, 250, 243, 253, 255, 255, 249, 214, 47, 18, 153, 130, 29, 32, 228, 245, 19, 8, 144, 126, 129, 127, 127, 140, 144, 143, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 139, 139, 138, 136, 148, 132, 151, 137, 252, 249, 140, 137, 251, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 252, 252, 252, 254, 255, 255, 255, 255, 255, 255, 250, 245, 238, 238, 255, 248, 255, 242, 231, 189, 0, 0, 79, 50, 59, 49, 61, 53, 53, 50, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 47, 49, 52, 51, 43, 42, 45, 49, 48, 54, 45, 45, 43, 42, 0, 0, 199, 185, 13, 0, 69, 97, 0, 26, 220, 235, 244, 254, 255, 255, 255, 248, 250, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 2, 2, 4, 0, 6, 0, 0, 0, 82, 78, 0, 0, 55, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 104, 101, 97, 106, 114, 0, 0, 139, 130, 132, 119, 118, 98, 104, 109, 100, 119, 113, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 113, 111, 111, 111, 115, 117, 122, 115, 106, 105, 122, 154, 126, 159, 0, 0, 138, 149, 118, 132, 0, 0, 116, 117, 132, 130, 104, 96, 105, 105, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 12, 20, 15, 12, 11, 18, 108, 122, 7, 12, 121, 126, 114, 115, 111, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 139, 138, 138, 139, 139, 139, 138, 138, 138, 138, 138, 139, 140, 141, 142, 142, 133, 131, 139, 6, 27, 214, 226, 247, 247, 255, 243, 251, 255, 244, 255, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 253, 251, 250, 252, 250, 246, 244, 253, 255, 215, 225, 16, 24, 211, 244, 240, 235, 24, 3, 134, 134, 146, 147, 130, 125, 134, 133, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 134, 142, 137, 134, 134, 143, 234, 252, 137, 144, 250, 255, 244, 251, 250, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 254, 248, 241, 241, 247, 245, 250, 232, 43, 0, 109, 67, 56, 38, 40, 26, 38, 51, 51, 68, 52, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 47, 45, 47, 52, 52, 45, 43, 45, 49, 58, 52, 35, 27, 38, 77, 61, 128, 0, 4, 122, 98, 45, 66, 0, 22, 220, 250, 255, 255, 255, 255, 252, 243, 252, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 5, 3, 0, 0, 0, 72, 82, 0, 0, 85, 81, 48, 45, 45, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 107, 107, 106, 106, 106, 106, 106, 106, 106, 107, 107, 108, 108, 107, 110, 107, 109, 104, 0, 0, 133, 126, 109, 109, 115, 108, 107, 114, 99, 116, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 111, 110, 110, 111, 115, 117, 117, 118, 117, 113, 116, 129, 125, 145, 0, 0, 126, 131, 115, 139, 0, 0, 121, 129, 109, 111, 114, 101, 114, 112, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 11, 19, 13, 14, 13, 15, 105, 112, 17, 19, 113, 117, 113, 115, 112, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 139, 139, 138, 137, 138, 138, 139, 139, 138, 138, 138, 137, 137, 137, 138, 139, 143, 139, 134, 136, 20, 33, 238, 247, 238, 246, 255, 255, 255, 255, 236, 249, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 253, 251, 250, 247, 250, 255, 253, 251, 254, 230, 234, 34, 44, 224, 250, 253, 252, 21, 3, 135, 146, 125, 131, 141, 132, 140, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 133, 141, 135, 136, 136, 140, 231, 242, 147, 151, 242, 248, 243, 251, 251, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 254, 252, 250, 255, 252, 250, 209, 6, 0, 75, 46, 32, 36, 44, 40, 43, 55, 45, 62, 52, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 47, 45, 47, 54, 54, 47, 43, 45, 47, 53, 55, 49, 40, 34, 48, 49, 92, 0, 0, 77, 64, 44, 84, 0, 20, 223, 254, 212, 218, 255, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 4, 1, 0, 0, 0, 69, 72, 0, 0, 77, 72, 47, 45, 46, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 106, 104, 104, 106, 106, 107, 107, 108, 110, 110, 111, 118, 107, 113, 106, 139, 131, 124, 112, 120, 124, 117, 115, 105, 118, 116, 130, 117, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 111, 108, 108, 111, 115, 117, 118, 117, 117, 114, 113, 114, 123, 128, 133, 106, 139, 105, 106, 122, 0, 0, 126, 106, 0, 0, 92, 111, 114, 108, 110, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 13, 17, 13, 13, 25, 7, 32, 16, 114, 107, 22, 16, 118, 115, 115, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 138, 138, 139, 140, 139, 139, 137, 137, 135, 135, 134, 134, 138, 128, 135, 148, 217, 238, 255, 253, 255, 254, 248, 249, 243, 255, 243, 255, 249, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 253, 254, 253, 251, 250, 248, 248, 255, 254, 252, 247, 246, 242, 240, 217, 255, 242, 250, 236, 21, 3, 141, 123, 12, 24, 123, 143, 140, 134, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 135, 139, 135, 135, 148, 132, 158, 146, 244, 239, 151, 147, 248, 251, 254, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 250, 255, 255, 255, 255, 255, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 247, 246, 198, 159, 96, 56, 34, 57, 66, 58, 54, 43, 55, 50, 63, 51, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 47, 45, 47, 54, 54, 49, 45, 43, 47, 54, 56, 55, 44, 35, 32, 42, 59, 85, 60, 77, 40, 54, 88, 0, 21, 222, 211, 56, 64, 203, 246, 255, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 2, 1, 0, 6, 0, 0, 0, 74, 68, 0, 0, 52, 45, 49, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 106, 104, 104, 106, 106, 107, 108, 110, 111, 111, 114, 117, 121, 124, 101, 142, 113, 111, 110, 115, 123, 112, 123, 110, 120, 118, 121, 117, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 110, 108, 108, 111, 115, 118, 117, 114, 115, 114, 115, 111, 122, 113, 111, 110, 113, 101, 116, 111, 0, 0, 114, 118, 0, 0, 112, 121, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 15, 18, 16, 3, 27, 12, 12, 11, 116, 115, 16, 10, 121, 114, 114, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 137, 138, 139, 140, 139, 139, 137, 136, 135, 134, 134, 134, 132, 138, 147, 150, 233, 236, 255, 255, 250, 250, 240, 254, 246, 255, 246, 248, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 253, 253, 251, 250, 247, 245, 253, 255, 255, 250, 255, 245, 242, 247, 255, 250, 255, 227, 35, 14, 144, 147, 13, 18, 146, 150, 132, 133, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 137, 140, 138, 125, 150, 137, 138, 141, 246, 247, 145, 141, 251, 250, 253, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 248, 250, 255, 255, 255, 255, 255, 252, 252, 252, 255, 255, 255, 255, 255, 255, 235, 226, 223, 165, 140, 67, 41, 38, 59, 72, 57, 64, 48, 55, 45, 47, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 47, 49, 56, 54, 51, 45, 43, 45, 51, 53, 56, 52, 44, 33, 41, 38, 50, 53, 48, 37, 66, 76, 0, 0, 182, 187, 2, 4, 183, 226, 243, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 4, 0, 8, 0, 0, 0, 76, 76, 0, 0, 55, 44, 48, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 107, 106, 104, 104, 104, 105, 106, 107, 107, 112, 107, 118, 116, 0, 0, 0, 0, 131, 120, 97, 111, 114, 118, 118, 115, 110, 108, 114, 115, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 110, 108, 110, 111, 115, 118, 118, 117, 113, 111, 110, 110, 113, 111, 107, 104, 101, 104, 114, 124, 135, 144, 0, 0, 148, 148, 0, 0, 110, 112, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 14, 18, 14, 23, 9, 12, 121, 118, 13, 14, 115, 123, 115, 117, 113, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 137, 138, 139, 139, 140, 138, 139, 137, 135, 136, 129, 140, 137, 0, 9, 8, 21, 229, 247, 244, 255, 249, 246, 248, 250, 254, 255, 253, 252, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 250, 252, 253, 253, 253, 252, 250, 248, 248, 250, 251, 253, 254, 254, 254, 254, 255, 255, 255, 251, 243, 231, 220, 25, 23, 217, 212, 13, 5, 136, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 136, 140, 136, 145, 132, 137, 247, 248, 143, 146, 244, 254, 245, 253, 252, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 250, 250, 255, 255, 255, 255, 255, 252, 251, 254, 255, 255, 255, 248, 252, 226, 46, 30, 23, 0, 108, 69, 32, 46, 59, 63, 54, 49, 45, 43, 40, 42, 47, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 52, 56, 54, 51, 45, 42, 43, 51, 56, 58, 54, 47, 42, 38, 40, 51, 52, 45, 43, 49, 67, 95, 130, 0, 0, 134, 134, 0, 50, 231, 255, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 3, 2, 8, 0, 0, 85, 78, 0, 0, 79, 78, 49, 47, 47, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 107, 106, 106, 104, 104, 104, 102, 106, 107, 106, 110, 118, 104, 120, 0, 0, 0, 0, 121, 124, 114, 111, 115, 117, 115, 113, 107, 107, 113, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 114, 110, 108, 110, 113, 117, 118, 118, 115, 113, 111, 110, 108, 108, 107, 104, 101, 101, 107, 118, 124, 121, 127, 0, 0, 130, 153, 0, 0, 120, 115, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 16, 20, 17, 13, 11, 17, 101, 113, 15, 22, 109, 116, 118, 116, 112, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 137, 138, 138, 139, 140, 140, 135, 137, 135, 132, 133, 142, 128, 149, 15, 28, 26, 61, 227, 253, 255, 253, 249, 248, 251, 253, 255, 255, 253, 252, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 250, 252, 253, 253, 252, 251, 250, 248, 249, 250, 251, 252, 254, 255, 255, 255, 255, 255, 255, 250, 246, 245, 237, 38, 39, 225, 235, 18, 5, 146, 142, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 138, 142, 139, 135, 134, 142, 227, 243, 145, 154, 238, 247, 248, 252, 251, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 252, 252, 255, 255, 255, 255, 254, 252, 250, 254, 255, 251, 245, 242, 214, 193, 0, 0, 0, 0, 75, 64, 50, 47, 56, 58, 47, 43, 43, 43, 42, 43, 47, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 52, 54, 56, 54, 49, 45, 42, 43, 51, 56, 59, 58, 52, 47, 40, 42, 47, 51, 49, 47, 43, 51, 63, 86, 0, 0, 83, 111, 0, 27, 231, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 1, 5, 5, 0, 0, 0, 65, 73, 0, 0, 73, 71, 52, 46, 46, 84, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 107, 106, 106, 104, 103, 104, 109, 109, 107, 114, 115, 106, 0, 0, 144, 144, 121, 111, 136, 118, 120, 118, 118, 117, 113, 110, 107, 110, 115, 117, 115, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 113, 110, 110, 111, 114, 117, 118, 117, 115, 113, 111, 110, 108, 107, 107, 107, 107, 107, 113, 124, 123, 108, 108, 128, 115, 137, 126, 0, 0, 106, 115, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 18, 17, 17, 12, 24, 9, 28, 17, 111, 110, 18, 16, 123, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 139, 140, 141, 140, 141, 139, 135, 139, 139, 129, 14, 14, 223, 240, 217, 216, 255, 244, 253, 251, 248, 250, 253, 255, 255, 252, 250, 249, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 251, 252, 252, 252, 252, 251, 250, 250, 249, 250, 250, 252, 253, 255, 255, 255, 255, 254, 251, 247, 248, 255, 253, 247, 226, 255, 221, 26, 19, 133, 145, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 140, 139, 139, 134, 147, 134, 154, 147, 241, 242, 147, 147, 253, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 254, 252, 254, 255, 255, 255, 255, 237, 205, 63, 4, 116, 88, 66, 54, 69, 46, 52, 50, 51, 49, 42, 40, 47, 52, 52, 52, 51, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 52, 54, 54, 52, 49, 45, 43, 43, 49, 54, 59, 59, 56, 52, 47, 45, 47, 49, 54, 51, 43, 40, 42, 52, 77, 61, 70, 67, 0, 27, 210, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 3, 2, 5, 0, 5, 0, 0, 0, 71, 71, 0, 0, 57, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 108, 106, 106, 104, 103, 103, 104, 108, 107, 111, 112, 118, 0, 0, 122, 138, 128, 134, 124, 109, 115, 117, 118, 115, 113, 111, 111, 114, 120, 120, 115, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 113, 110, 110, 113, 115, 118, 118, 115, 114, 113, 111, 111, 110, 108, 108, 110, 111, 113, 117, 124, 120, 103, 101, 113, 128, 125, 127, 0, 0, 101, 114, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 16, 14, 25, 7, 25, 7, 122, 117, 11, 6, 121, 116, 116, 128, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 137, 138, 139, 140, 141, 140, 139, 137, 135, 137, 135, 142, 4, 19, 223, 255, 252, 255, 253, 238, 243, 245, 249, 252, 254, 254, 252, 250, 247, 247, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 250, 251, 252, 253, 252, 251, 250, 250, 251, 251, 250, 251, 251, 252, 253, 254, 254, 253, 250, 248, 247, 250, 255, 255, 252, 254, 248, 223, 22, 8, 128, 146, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 139, 139, 138, 136, 148, 132, 151, 137, 252, 249, 140, 137, 251, 252, 255, 237, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 252, 250, 254, 255, 255, 255, 250, 228, 206, 37, 0, 85, 67, 54, 58, 47, 34, 46, 48, 47, 42, 38, 40, 49, 54, 56, 56, 51, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 52, 52, 52, 51, 49, 45, 43, 45, 47, 51, 56, 58, 58, 54, 51, 47, 43, 47, 56, 56, 45, 38, 38, 40, 47, 56, 53, 72, 0, 21, 207, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 2, 2, 4, 0, 6, 0, 0, 0, 82, 78, 0, 0, 55, 46, 50, 82, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 108, 108, 106, 106, 104, 103, 103, 104, 107, 109, 113, 114, 120, 0, 0, 131, 118, 97, 102, 115, 122, 121, 123, 117, 115, 114, 115, 118, 121, 124, 123, 117, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 113, 111, 110, 110, 114, 117, 120, 118, 115, 113, 111, 111, 113, 111, 110, 110, 114, 115, 118, 120, 120, 115, 104, 101, 107, 102, 127, 156, 0, 0, 127, 102, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 12, 20, 15, 12, 11, 18, 108, 122, 7, 12, 121, 126, 114, 115, 111, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 137, 136, 138, 138, 140, 141, 140, 139, 139, 134, 136, 134, 140, 3, 18, 235, 252, 239, 245, 255, 255, 249, 251, 251, 252, 253, 251, 249, 247, 245, 246, 249, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 253, 251, 250, 249, 250, 251, 252, 252, 252, 251, 251, 252, 253, 253, 252, 247, 246, 248, 251, 255, 255, 251, 233, 239, 236, 15, 3, 157, 135, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 134, 142, 137, 134, 134, 143, 234, 252, 137, 144, 250, 255, 244, 251, 250, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 254, 252, 254, 255, 255, 255, 252, 229, 209, 41, 0, 112, 69, 33, 29, 45, 54, 52, 54, 43, 40, 40, 43, 49, 51, 52, 52, 51, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 51, 51, 49, 47, 47, 45, 45, 45, 45, 47, 51, 52, 54, 54, 52, 47, 40, 42, 56, 58, 51, 47, 51, 49, 40, 33, 69, 123, 0, 37, 245, 250, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 5, 3, 0, 0, 0, 72, 82, 0, 0, 85, 81, 48, 45, 45, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 110, 108, 106, 104, 103, 101, 101, 107, 108, 109, 116, 118, 109, 0, 0, 133, 110, 130, 109, 110, 110, 107, 116, 115, 114, 115, 117, 121, 123, 123, 120, 117, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 113, 111, 110, 111, 115, 118, 120, 118, 114, 111, 111, 111, 114, 114, 111, 113, 114, 117, 121, 120, 115, 111, 108, 108, 103, 139, 136, 137, 0, 0, 96, 108, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 11, 19, 13, 14, 13, 15, 105, 112, 17, 19, 113, 117, 113, 115, 112, 131, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 136, 136, 137, 138, 140, 141, 141, 142, 140, 134, 138, 137, 127, 11, 12, 218, 229, 255, 253, 253, 249, 239, 247, 252, 253, 251, 250, 248, 247, 247, 248, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 252, 254, 253, 251, 250, 248, 249, 252, 253, 253, 253, 251, 250, 252, 252, 252, 250, 246, 247, 251, 253, 252, 253, 247, 255, 229, 198, 25, 0, 128, 143, 138, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 133, 141, 135, 136, 136, 140, 231, 242, 147, 151, 242, 248, 243, 251, 251, 240, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 252, 252, 255, 255, 255, 255, 240, 211, 70, 14, 133, 77, 73, 41, 47, 46, 42, 45, 38, 36, 43, 45, 47, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 45, 43, 45, 45, 47, 47, 43, 43, 45, 47, 51, 52, 52, 49, 43, 45, 56, 56, 47, 45, 56, 54, 36, 77, 97, 131, 33, 62, 227, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 4, 1, 0, 0, 0, 69, 72, 0, 0, 77, 72, 47, 45, 46, 85, 0, 28, 228, 255, 254, 255, 255, 255, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 110, 110, 108, 106, 104, 103, 101, 101, 100, 105, 109, 109, 114, 125, 113, 124, 0, 0, 117, 116, 112, 105, 114, 119, 111, 111, 114, 117, 120, 118, 114, 111, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 113, 111, 110, 111, 115, 118, 120, 118, 113, 110, 110, 111, 114, 115, 114, 113, 113, 115, 121, 118, 108, 108, 117, 120, 124, 111, 0, 0, 109, 116, 112, 93, 106, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 121, 0, 0, 133, 111, 118, 116, 115, 110, 14, 11, 13, 16, 113, 116, 114, 114, 114, 114, 114, 114, 114, 114, 12, 15, 113, 116, 116, 113, 15, 12, 16, 16, 16, 16, 16, 16, 16, 16, 13, 17, 13, 13, 25, 7, 32, 16, 114, 107, 22, 16, 118, 115, 115, 130, 0, 0, 118, 108, 102, 105, 105, 111, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 136, 135, 136, 137, 139, 141, 142, 136, 138, 135, 130, 130, 137, 123, 146, 17, 50, 227, 247, 252, 247, 252, 255, 255, 255, 252, 250, 248, 250, 251, 252, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 253, 254, 254, 251, 249, 248, 249, 253, 255, 255, 254, 251, 250, 250, 251, 251, 249, 246, 249, 255, 255, 249, 246, 255, 226, 30, 18, 130, 139, 148, 132, 139, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 135, 142, 0, 17, 237, 247, 250, 252, 254, 249, 145, 139, 138, 143, 247, 253, 251, 251, 251, 251, 251, 251, 251, 248, 141, 144, 247, 253, 253, 247, 144, 138, 139, 139, 138, 138, 138, 138, 138, 139, 135, 139, 135, 135, 148, 132, 158, 146, 244, 239, 151, 147, 248, 251, 254, 239, 19, 0, 142, 139, 139, 142, 133, 137, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 252, 255, 255, 255, 255, 255, 254, 250, 248, 253, 255, 255, 251, 249, 220, 196, 0, 0, 66, 55, 57, 49, 52, 48, 35, 35, 45, 49, 47, 45, 47, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 45, 42, 42, 43, 47, 49, 47, 43, 40, 40, 42, 47, 49, 52, 52, 54, 54, 56, 49, 35, 35, 54, 58, 58, 61, 0, 11, 187, 233, 255, 249, 255, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 233, 30, 0, 90, 49, 52, 48, 49, 58, 0, 2, 2, 0, 64, 53, 49, 47, 49, 49, 51, 51, 51, 63, 0, 0, 62, 51, 53, 64, 0, 2, 0, 0, 1, 3, 3, 1, 1, 0, 0, 2, 1, 0, 6, 0, 0, 0, 74, 68, 0, 0, 52, 45, 49, 84, 0, 28, 228, 255, 254, 255, 255, 255, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 127, 121, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 132, 131, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 127, 121, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 132, 131, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 127, 121, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 134, 132, 131, 129, 127, 125, 125, 124, 124, 124, 127, 129, 131, 137, 132, 145, 138, 0, 0, 168, 158, 140, 134, 154, 143, 142, 142, 142, 144, 146, 146, 144, 144, 144, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 142, 135, 137, 144, 146, 144, 145, 149, 149, 145, 142, 139, 141, 144, 146, 148, 148, 144, 145, 149, 148, 138, 139, 151, 153, 149, 157, 0, 0, 149, 139, 119, 123, 120, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 132, 131, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 127, 121, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 132, 131, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 127, 121, 122, 131, 132, 127, 127, 129, 131, 131, 129, 127, 127, 128, 129, 132, 132, 130, 139, 4, 0, 160, 142, 147, 146, 146, 141, 45, 42, 43, 46, 144, 144, 137, 138, 146, 148, 142, 142, 145, 146, 44, 46, 141, 144, 146, 144, 49, 47, 47, 45, 45, 45, 45, 45, 45, 45, 44, 47, 45, 32, 56, 41, 41, 40, 139, 139, 49, 44, 148, 143, 145, 159, 0, 4, 135, 126, 123, 127, 129, 136, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 134, 134, 134, 133, 134, 134, 135, 138, 138, 136, 136, 134, 131, 131, 124, 134, 135, 9, 17, 224, 233, 231, 229, 245, 233, 236, 235, 233, 232, 231, 232, 234, 234, 233, 231, 231, 231, 231, 231, 231, 231, 231, 231, 231, 231, 231, 231, 231, 232, 235, 235, 234, 233, 233, 231, 229, 230, 233, 235, 235, 235, 233, 231, 231, 230, 231, 230, 228, 230, 238, 237, 228, 225, 230, 221, 16, 0, 147, 139, 130, 142, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 138, 138, 135, 135, 136, 136, 135, 135, 135, 135, 136, 136, 136, 136, 135, 135, 133, 139, 0, 10, 221, 227, 231, 232, 234, 230, 127, 122, 121, 126, 228, 234, 234, 234, 232, 231, 232, 232, 231, 229, 123, 127, 230, 234, 234, 229, 126, 120, 122, 122, 122, 122, 122, 122, 122, 122, 121, 124, 121, 109, 133, 120, 121, 123, 231, 231, 128, 122, 233, 231, 234, 224, 11, 0, 140, 138, 137, 139, 131, 134, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 206, 209, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 206, 209, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 204, 208, 213, 220, 224, 225, 220, 213, 209, 208, 211, 216, 217, 219, 209, 212, 182, 4, 0, 99, 78, 78, 73, 80, 60, 54, 56, 68, 72, 67, 61, 59, 61, 67, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 72, 75, 72, 58, 56, 67, 70, 68, 65, 61, 59, 63, 63, 65, 65, 63, 67, 75, 77, 75, 67, 54, 56, 74, 79, 73, 98, 0, 9, 197, 213, 209, 221, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 206, 209, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 206, 209, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 220, 216, 206, 204, 213, 215, 209, 208, 208, 209, 213, 213, 211, 208, 204, 206, 212, 199, 9, 0, 100, 71, 73, 71, 70, 78, 1, 9, 9, 3, 81, 76, 77, 74, 63, 63, 72, 74, 68, 77, 0, 0, 80, 74, 72, 76, 0, 2, 4, 6, 10, 10, 10, 10, 8, 8, 7, 12, 12, 0, 17, 0, 0, 0, 98, 96, 0, 0, 77, 67, 68, 94, 0, 5, 195, 214, 210, 211, 205, 207, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 229, 6, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 229, 6, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 229, 6, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 237, 236, 236, 235, 235, 235, 235, 235, 236, 236, 237, 239, 239, 240, 233, 10, 14, 118, 110, 223, 219, 219, 237, 229, 229, 219, 220, 114, 114, 116, 113, 229, 226, 226, 226, 226, 226, 226, 226, 226, 226, 226, 226, 226, 226, 226, 219, 0, 3, 111, 108, 225, 222, 221, 239, 229, 229, 219, 218, 113, 114, 117, 114, 229, 226, 228, 228, 225, 225, 229, 229, 228, 230, 237, 240, 239, 237, 235, 226, 4, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 229, 6, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 236, 229, 6, 14, 123, 119, 234, 231, 229, 247, 240, 239, 228, 228, 123, 123, 127, 125, 240, 239, 242, 239, 230, 226, 228, 226, 226, 226, 226, 226, 226, 226, 226, 219, 0, 4, 113, 109, 225, 221, 219, 237, 230, 229, 219, 218, 113, 114, 117, 115, 230, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 219, 0, 4, 113, 109, 226, 221, 219, 242, 243, 245, 231, 228, 121, 122, 127, 128, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 198, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 198, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 198, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 195, 195, 195, 196, 196, 197, 197, 197, 196, 196, 195, 194, 194, 194, 198, 0, 7, 90, 84, 220, 220, 208, 221, 215, 218, 214, 214, 107, 102, 95, 91, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 215, 12, 17, 96, 87, 220, 219, 207, 220, 214, 218, 214, 216, 108, 101, 94, 90, 213, 213, 212, 213, 215, 215, 211, 211, 212, 209, 202, 198, 196, 196, 196, 199, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 198, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 198, 0, 0, 78, 69, 203, 202, 191, 203, 196, 201, 197, 198, 90, 84, 77, 73, 195, 196, 197, 202, 209, 213, 212, 213, 213, 212, 211, 210, 210, 211, 212, 215, 12, 16, 95, 86, 220, 219, 208, 220, 211, 215, 213, 215, 107, 101, 92, 87, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 211, 214, 11, 15, 94, 85, 219, 219, 208, 217, 202, 202, 197, 198, 91, 85, 77, 72, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 203, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 189, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 203, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 189, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 203, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 189, 196, 199, 199, 201, 199, 196, 196, 196, 196, 197, 197, 197, 197, 194, 192, 0, 0, 6, 0, 141, 144, 119, 126, 118, 126, 133, 136, 19, 4, 0, 0, 126, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 141, 0, 0, 0, 0, 136, 142, 119, 128, 119, 126, 132, 133, 17, 5, 0, 0, 128, 135, 135, 132, 128, 128, 135, 137, 134, 142, 160, 176, 187, 194, 197, 204, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 189, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 203, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 189, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 203, 9, 4, 59, 46, 200, 204, 182, 190, 183, 192, 195, 198, 81, 67, 54, 52, 190, 190, 176, 160, 142, 135, 134, 134, 134, 137, 144, 148, 148, 144, 137, 141, 0, 0, 0, 0, 138, 142, 119, 132, 132, 140, 137, 136, 19, 9, 0, 3, 139, 146, 148, 148, 148, 148, 146, 146, 146, 148, 148, 148, 146, 144, 141, 148, 0, 0, 2, 0, 139, 142, 119, 137, 148, 170, 188, 198, 81, 69, 54, 45, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 149, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 249, 26, 20, 151, 168, 235, 255, 255, 255, 255, 255, 255, 254, 129, 111, 155, 152, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 197, 5, 0, 89, 94, 179, 201, 198, 188, 188, 201, 202, 201, 82, 59, 86, 77, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 18, 142, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 160, 0, 0, 32, 31, 132, 155, 141, 123, 125, 142, 155, 157, 38, 11, 27, 12, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 143, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 131, 16, 18, 241, 240, 159, 142, 156, 159, 158, 156, 143, 132, 29, 48, 222, 255, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 201, 74, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 77, 0, 4, 192, 175, 94, 72, 77, 74, 73, 77, 68, 72, 0, 14, 172, 202, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 154, 15, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 31, 0, 0, 152, 121, 38, 10, 2, 0, 0, 2, 1, 20, 0, 0, 135, 159, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 150, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 156, 157, 141, 15, 11, 254, 255, 140, 145, 160, 165, 157, 164, 159, 147, 25, 24, 240, 255, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 206, 79, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 78, 77, 81, 0, 0, 210, 202, 70, 67, 75, 76, 71, 79, 76, 82, 0, 2, 198, 207, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 162, 15, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 3, 4, 27, 0, 0, 181, 153, 8, 0, 0, 0, 0, 0, 0, 24, 0, 0, 173, 173, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 251, 150, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 155, 157, 141, 36, 20, 240, 254, 143, 161, 153, 150, 157, 161, 160, 147, 22, 15, 242, 246, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 187, 73, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 72, 71, 75, 4, 0, 193, 192, 68, 82, 74, 71, 75, 78, 71, 77, 0, 0, 197, 188, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 139, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 165, 145, 1, 5, 0, 0, 0, 0, 0, 15, 0, 0, 168, 150, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 252, 153, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 145, 27, 21, 250, 255, 146, 155, 147, 159, 157, 160, 159, 148, 23, 14, 245, 245, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 188, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 77, 0, 0, 205, 201, 71, 73, 68, 77, 75, 75, 67, 77, 0, 0, 201, 190, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 140, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 176, 157, 4, 0, 0, 3, 0, 0, 0, 13, 0, 0, 172, 151, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 255, 150, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 141, 26, 15, 240, 253, 141, 150, 160, 161, 164, 166, 164, 152, 27, 22, 239, 247, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 199, 76, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 79, 0, 0, 196, 192, 70, 70, 74, 71, 71, 71, 69, 78, 0, 4, 202, 201, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 154, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 0, 0, 167, 147, 8, 0, 0, 0, 0, 0, 0, 15, 0, 0, 176, 167, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 255, 145, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 136, 22, 13, 245, 255, 138, 140, 160, 150, 160, 161, 156, 142, 27, 23, 229, 248, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 202, 74, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 73, 72, 77, 0, 0, 202, 201, 75, 70, 81, 64, 70, 71, 68, 73, 0, 0, 192, 203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 160, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 170, 157, 24, 11, 14, 0, 0, 0, 0, 16, 0, 0, 165, 170, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 255, 146, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 151, 152, 135, 17, 16, 243, 255, 36, 36, 140, 145, 150, 149, 139, 132, 29, 31, 237, 252, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 201, 75, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 75, 74, 79, 0, 0, 195, 196, 0, 0, 80, 77, 76, 75, 70, 75, 0, 0, 192, 202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 156, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 159, 152, 0, 0, 28, 16, 11, 12, 15, 30, 0, 0, 161, 169, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 255, 148, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 137, 18, 29, 245, 244, 40, 27, 115, 131, 132, 124, 134, 118, 42, 37, 252, 254, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 75, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 78, 0, 10, 192, 187, 9, 1, 77, 82, 78, 72, 86, 75, 3, 0, 196, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 144, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 150, 142, 0, 0, 41, 39, 31, 25, 50, 43, 0, 0, 159, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 153, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 141, 30, 21, 148, 134, 14, 4, 22, 21, 24, 32, 21, 24, 119, 118, 255, 255, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 90, 80, 0, 0, 4, 0, 0, 2, 0, 0, 80, 69, 202, 191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 133, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 49, 28, 154, 138, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 155, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 156, 158, 142, 25, 20, 153, 127, 27, 7, 15, 21, 22, 35, 21, 32, 112, 124, 255, 255, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 75, 0, 0, 96, 73, 5, 0, 0, 0, 0, 7, 0, 3, 77, 76, 197, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 49, 38, 149, 139, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 255, 152, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 158, 159, 141, 15, 28, 229, 255, 227, 240, 242, 255, 250, 244, 249, 231, 37, 32, 246, 252, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 192, 73, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 75, 0, 15, 183, 205, 189, 205, 197, 208, 198, 194, 204, 194, 9, 0, 196, 193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 142, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 7, 147, 163, 166, 185, 166, 171, 161, 159, 175, 168, 0, 0, 159, 149, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 152, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 139, 14, 10, 229, 255, 247, 255, 255, 255, 255, 255, 255, 249, 21, 20, 243, 255, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 205, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 76, 0, 0, 188, 210, 192, 209, 196, 192, 194, 192, 202, 201, 0, 0, 198, 207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 159, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 160, 170, 153, 166, 146, 139, 142, 142, 155, 165, 0, 0, 167, 168, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 255, 152, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 141, 20, 16, 252, 246, 152, 140, 152, 157, 148, 158, 143, 141, 21, 32, 231, 254, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 76, 0, 0, 206, 181, 77, 61, 72, 78, 70, 80, 65, 79, 0, 7, 180, 190, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 143, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 182, 139, 19, 0, 3, 11, 4, 14, 0, 30, 0, 2, 153, 152, 156, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 152, 155, 153, 153, 155, 156, 155, 155, 155, 155, 158, 156, 153, 153, 155, 141, 28, 17, 247, 252, 164, 162, 167, 148, 154, 152, 164, 139, 21, 17, 244, 255, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 74, 74, 74, 74, 74, 73, 73, 74, 74, 74, 73, 74, 74, 74, 74, 76, 0, 0, 201, 185, 80, 71, 81, 66, 72, 70, 80, 74, 0, 0, 193, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 144, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 177, 140, 10, 0, 6, 0, 0, 0, 7, 20, 0, 0, 164, 155, 162, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 158, 155, 144, 159, 151, 166, 158, 151, 159, 159, 159, 159, 157, 146, 164, 138, 21, 22, 237, 253, 157, 151, 152, 150, 151, 156, 159, 135, 19, 14, 245, 255, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 204, 76, 73, 70, 84, 67, 80, 75, 71, 77, 77, 70, 73, 81, 72, 80, 72, 0, 4, 198, 191, 73, 60, 73, 73, 69, 73, 79, 73, 0, 0, 195, 205, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 148, 0, 0, 0, 16, 0, 7, 5, 0, 1, 0, 0, 0, 6, 1, 8, 14, 0, 0, 167, 140, 0, 0, 4, 5, 0, 0, 8, 22, 0, 0, 162, 159, 155, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 248, 150, 163, 147, 158, 156, 153, 155, 148, 151, 157, 161, 159, 154, 144, 160, 141, 23, 11, 237, 255, 153, 161, 154, 144, 159, 159, 141, 139, 17, 15, 246, 244, 72, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 73, 81, 70, 79, 67, 62, 72, 68, 69, 75, 73, 75, 78, 70, 78, 76, 0, 0, 202, 199, 71, 71, 79, 71, 76, 72, 61, 79, 0, 0, 200, 183, 0, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 129, 1, 5, 2, 12, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 5, 20, 0, 0, 172, 149, 0, 0, 12, 3, 0, 0, 0, 27, 0, 0, 166, 138, 151, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 147, 156, 151, 159, 174, 164, 167, 154, 155, 160, 158, 152, 149, 145, 150, 140, 21, 8, 231, 254, 144, 158, 154, 147, 155, 165, 145, 146, 17, 11, 247, 255, 79, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 201, 80, 78, 64, 66, 79, 72, 82, 71, 73, 79, 77, 74, 72, 69, 72, 81, 2, 0, 201, 201, 66, 72, 79, 72, 68, 74, 61, 85, 0, 0, 206, 202, 20, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 155, 25, 16, 0, 0, 11, 5, 15, 3, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 177, 157, 0, 0, 12, 4, 0, 0, 0, 31, 0, 0, 174, 160, 139, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 240, 135, 129, 161, 154, 157, 154, 157, 154, 156, 159, 157, 158, 159, 157, 132, 124, 20, 45, 219, 253, 163, 152, 147, 151, 166, 168, 150, 138, 14, 25, 210, 238, 80, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 194, 82, 63, 77, 61, 68, 67, 70, 66, 69, 72, 74, 77, 80, 83, 71, 77, 0, 24, 180, 195, 83, 66, 70, 73, 75, 75, 66, 78, 0, 16, 180, 195, 38, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 160, 42, 13, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 10, 6, 31, 0, 5, 147, 147, 14, 0, 0, 1, 0, 0, 0, 26, 0, 9, 156, 163, 31, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 24, 28, 41, 145, 154, 146, 153, 163, 179, 172, 169, 163, 159, 152, 130, 47, 26, 249, 220, 157, 151, 149, 161, 163, 153, 165, 156, 157, 130, 19, 0, 33, 21, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 75, 75, 70, 73, 72, 82, 72, 70, 70, 72, 68, 62, 9, 0, 211, 172, 96, 76, 58, 69, 81, 71, 72, 63, 74, 74, 5, 0, 15, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 0, 0, 23, 16, 12, 10, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 175, 126, 42, 11, 0, 0, 7, 0, 0, 0, 4, 27, 0, 2, 5, 0, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 22, 43, 113, 143, 139, 140, 153, 154, 165, 162, 159, 159, 158, 138, 27, 14, 239, 255, 146, 151, 167, 154, 154, 154, 157, 154, 167, 130, 22, 4, 22, 22, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 8, 61, 82, 81, 73, 73, 62, 70, 67, 69, 76, 78, 79, 7, 0, 192, 198, 75, 71, 76, 63, 72, 72, 64, 61, 84, 72, 4, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 21, 35, 33, 20, 4, 0, 0, 0, 0, 0, 5, 23, 0, 0, 148, 138, 11, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 233, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 254, 237, 201, 49, 28, 29, 40, 142, 155, 150, 149, 147, 146, 143, 128, 14, 11, 245, 255, 144, 149, 155, 147, 148, 152, 164, 166, 165, 132, 30, 36, 222, 255, 206, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 205, 173, 15, 0, 0, 0, 79, 84, 80, 77, 78, 79, 76, 82, 5, 2, 195, 201, 73, 72, 73, 65, 74, 75, 74, 73, 78, 66, 0, 14, 184, 212, 187, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 187, 184, 151, 0, 0, 0, 0, 25, 18, 10, 3, 1, 1, 0, 20, 0, 0, 146, 139, 9, 4, 0, 0, 3, 3, 0, 0, 7, 14, 0, 1, 161, 183, 240, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 240, 243, 246, 25, 22, 41, 29, 134, 118, 123, 125, 131, 133, 125, 119, 14, 25, 255, 255, 149, 155, 148, 154, 150, 147, 154, 160, 150, 143, 29, 22, 247, 241, 202, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 200, 210, 0, 0, 9, 0, 89, 70, 77, 79, 85, 84, 76, 81, 0, 2, 196, 186, 75, 80, 70, 77, 80, 72, 67, 70, 66, 76, 0, 0, 203, 191, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 166, 176, 0, 0, 0, 0, 48, 22, 27, 27, 26, 25, 17, 32, 0, 0, 142, 121, 10, 13, 0, 5, 11, 4, 0, 0, 0, 23, 0, 0, 176, 158, 149, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 243, 145, 124, 253, 228, 237, 245, 25, 20, 19, 22, 17, 20, 25, 28, 241, 250, 146, 153, 151, 151, 152, 151, 148, 151, 158, 156, 151, 141, 31, 21, 244, 239, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 86, 69, 209, 190, 198, 208, 0, 0, 0, 5, 0, 0, 0, 0, 203, 197, 73, 73, 73, 74, 73, 74, 75, 74, 72, 70, 73, 81, 0, 0, 207, 194, 17, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 154, 28, 5, 162, 153, 165, 181, 0, 0, 0, 0, 0, 0, 0, 0, 184, 166, 18, 4, 7, 6, 4, 2, 7, 4, 0, 0, 7, 31, 0, 0, 181, 165, 150, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 247, 142, 152, 255, 255, 251, 219, 50, 20, 17, 14, 14, 27, 11, 23, 251, 254, 154, 157, 154, 154, 155, 155, 154, 155, 160, 151, 153, 139, 29, 22, 240, 239, 68, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 194, 70, 79, 193, 207, 196, 170, 14, 0, 0, 0, 0, 10, 0, 0, 200, 186, 74, 75, 76, 76, 75, 76, 76, 75, 74, 67, 79, 80, 0, 0, 202, 195, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 154, 0, 0, 132, 160, 155, 138, 0, 0, 0, 0, 0, 0, 0, 0, 183, 151, 13, 2, 4, 4, 2, 1, 4, 2, 0, 0, 18, 36, 0, 0, 181, 170, 176, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 255, 165, 161, 160, 148, 141, 168, 231, 255, 240, 251, 249, 212, 27, 13, 239, 255, 150, 152, 151, 152, 155, 157, 158, 160, 169, 154, 149, 131, 29, 26, 244, 246, 80, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 196, 82, 70, 77, 67, 59, 93, 172, 206, 190, 206, 210, 187, 17, 0, 189, 195, 73, 73, 74, 73, 72, 72, 71, 71, 78, 68, 74, 72, 0, 0, 201, 198, 0, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 159, 12, 0, 9, 11, 9, 51, 138, 175, 153, 167, 177, 165, 15, 0, 166, 151, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 0, 0, 182, 176, 150, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 249, 141, 161, 155, 157, 151, 155, 254, 255, 255, 255, 248, 222, 23, 20, 244, 255, 148, 152, 151, 152, 155, 157, 158, 158, 154, 152, 125, 124, 45, 34, 251, 241, 60, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 189, 61, 72, 69, 72, 62, 73, 182, 200, 200, 195, 195, 186, 9, 2, 194, 190, 73, 73, 74, 73, 72, 72, 71, 71, 68, 73, 61, 74, 8, 0, 205, 190, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 153, 0, 0, 0, 7, 2, 17, 132, 151, 142, 137, 145, 150, 0, 0, 169, 145, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 41, 0, 0, 189, 171, 144, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 255, 139, 150, 149, 150, 155, 136, 160, 148, 158, 149, 146, 144, 25, 25, 241, 255, 149, 154, 153, 153, 153, 153, 154, 152, 150, 137, 46, 35, 20, 21, 245, 250, 79, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 203, 78, 83, 80, 78, 80, 59, 85, 69, 75, 70, 78, 94, 0, 0, 197, 201, 76, 75, 75, 75, 75, 75, 75, 75, 80, 77, 2, 3, 0, 0, 202, 202, 0, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 166, 11, 4, 3, 6, 12, 0, 18, 0, 0, 0, 15, 45, 0, 0, 170, 159, 8, 0, 0, 0, 0, 0, 0, 5, 18, 25, 0, 0, 0, 0, 185, 180, 126, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 246, 129, 125, 129, 124, 139, 140, 136, 141, 133, 139, 135, 122, 47, 51, 234, 255, 140, 141, 139, 137, 137, 137, 137, 134, 128, 117, 21, 17, 32, 48, 236, 249, 86, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 192, 84, 83, 82, 75, 88, 85, 75, 77, 67, 77, 79, 74, 2, 5, 184, 201, 78, 78, 79, 80, 80, 80, 80, 81, 81, 79, 0, 0, 9, 16, 186, 190, 27, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 148, 29, 25, 26, 19, 35, 31, 18, 16, 7, 18, 28, 28, 0, 0, 151, 162, 27, 24, 25, 27, 25, 25, 25, 29, 35, 42, 0, 0, 0, 0, 153, 150, 14, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 143, 27, 14, 17, 15, 14, 15, 21, 23, 27, 18, 14, 31, 120, 143, 255, 252, 29, 21, 18, 17, 15, 15, 18, 17, 14, 24, 8, 25, 101, 101, 161, 156, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 77, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 61, 73, 204, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 13, 76, 57, 92, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 159, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 10, 27, 0, 5, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 144, 23, 8, 3, 6, 0, 8, 7, 7, 0, 0, 0, 18, 150, 150, 255, 250, 21, 7, 3, 1, 0, 1, 3, 3, 4, 5, 1, 8, 116, 138, 145, 163, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 74, 0, 3, 0, 3, 0, 5, 0, 1, 1, 7, 0, 0, 86, 68, 185, 194, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 1, 88, 88, 67, 70, 6, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 0, 9, 4, 10, 7, 12, 0, 3, 14, 21, 9, 0, 42, 10, 133, 159, 0, 5, 9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 0
);


begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   blue <= std_logic_vector(to_unsigned(ROM(addr_reg),8));
	
end arch;

